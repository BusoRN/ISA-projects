library verilog;
use verilog.vl_types.all;
entity tb_acs4 is
end tb_acs4;
