
module FIR ( DIN, H0, H1, H2, H3, H4, H5, H6, VIN, RST_n, CLK, VOUT, DOUT );
  input [7:0] DIN;
  input [7:0] H0;
  input [7:0] H1;
  input [7:0] H2;
  input [7:0] H3;
  input [7:0] H4;
  input [7:0] H5;
  input [7:0] H6;
  output [7:0] DOUT;
  input VIN, RST_n, CLK;
  output VOUT;
  wire   SR_to_MUX, MUX_to_PIPE1, PIPE1_to_PIPE2, PIPE2_to_REGOUT,
         ADD_esteso_0__17_, ADD_esteso_0__14_, ADD_esteso_0__13_,
         ADD_esteso_0__12_, ADD_esteso_0__11_, ADD_esteso_0__10_,
         ADD_esteso_0__9_, ADD_esteso_0__8_, ADD_esteso_0__7_,
         ADD_esteso_0__6_, ADD_esteso_0__5_, ADD_esteso_0__4_,
         ADD_esteso_0__3_, ADD_esteso_0__2_, ADD_esteso_0__1_,
         ADD_esteso_0__0_, ADD_esteso_1__17_, ADD_esteso_1__14_,
         ADD_esteso_1__13_, ADD_esteso_1__12_, ADD_esteso_1__11_,
         ADD_esteso_1__10_, ADD_esteso_1__9_, ADD_esteso_1__8_,
         ADD_esteso_1__7_, ADD_esteso_1__6_, ADD_esteso_1__5_,
         ADD_esteso_1__4_, ADD_esteso_1__3_, ADD_esteso_1__2_,
         ADD_esteso_1__1_, ADD_esteso_1__0_, ADD_esteso_2__17_,
         ADD_esteso_2__14_, ADD_esteso_2__13_, ADD_esteso_2__12_,
         ADD_esteso_2__11_, ADD_esteso_2__10_, ADD_esteso_2__9_,
         ADD_esteso_2__8_, ADD_esteso_2__7_, ADD_esteso_2__6_,
         ADD_esteso_2__5_, ADD_esteso_2__4_, ADD_esteso_2__3_,
         ADD_esteso_2__2_, ADD_esteso_2__1_, ADD_esteso_2__0_,
         ADD_esteso_3__17_, ADD_esteso_3__14_, ADD_esteso_3__13_,
         ADD_esteso_3__12_, ADD_esteso_3__11_, ADD_esteso_3__10_,
         ADD_esteso_3__9_, ADD_esteso_3__8_, ADD_esteso_3__7_,
         ADD_esteso_3__6_, ADD_esteso_3__5_, ADD_esteso_3__4_,
         ADD_esteso_3__3_, ADD_esteso_3__2_, ADD_esteso_3__1_,
         ADD_esteso_3__0_, ADD_esteso_4__17_, ADD_esteso_4__14_,
         ADD_esteso_4__13_, ADD_esteso_4__12_, ADD_esteso_4__11_,
         ADD_esteso_4__10_, ADD_esteso_4__9_, ADD_esteso_4__8_,
         ADD_esteso_4__7_, ADD_esteso_4__6_, ADD_esteso_4__5_,
         ADD_esteso_4__4_, ADD_esteso_4__3_, ADD_esteso_4__2_,
         ADD_esteso_4__1_, ADD_esteso_4__0_, ADD_esteso_5__17_,
         ADD_esteso_5__14_, ADD_esteso_5__13_, ADD_esteso_5__12_,
         ADD_esteso_5__11_, ADD_esteso_5__10_, ADD_esteso_5__9_,
         ADD_esteso_5__8_, ADD_esteso_5__7_, ADD_esteso_5__6_,
         ADD_esteso_5__5_, ADD_esteso_5__4_, ADD_esteso_5__3_,
         ADD_esteso_5__2_, ADD_esteso_5__1_, ADD_esteso_5__0_,
         ADD_esteso_6__17_, ADD_esteso_6__14_, ADD_esteso_6__13_,
         ADD_esteso_6__12_, ADD_esteso_6__11_, ADD_esteso_6__10_,
         ADD_esteso_6__9_, ADD_esteso_6__8_, ADD_esteso_6__7_,
         ADD_esteso_6__6_, ADD_esteso_6__5_, ADD_esteso_6__4_,
         ADD_esteso_6__3_, ADD_esteso_6__2_, ADD_esteso_6__1_,
         ADD_esteso_6__0_, ADD_esteso_10__17_, ADD_esteso_10__16_,
         ADD_esteso_10__15_, ADD_esteso_10__14_, ADD_esteso_10__13_,
         ADD_esteso_10__12_, ADD_esteso_10__11_, ADD_esteso_10__10_,
         ADD_esteso_10__9_, ADD_esteso_10__8_, ADD_esteso_10__7_,
         ADD_esteso_10__6_, ADD_esteso_10__5_, ADD_esteso_10__4_,
         ADD_esteso_10__3_, ADD_esteso_10__2_, ADD_esteso_10__1_,
         ADD_esteso_10__0_, ADD_esteso_11__17_, ADD_esteso_11__16_,
         ADD_esteso_11__15_, ADD_esteso_11__14_, ADD_esteso_11__13_,
         ADD_esteso_11__12_, ADD_esteso_11__11_, ADD_esteso_11__10_,
         ADD_esteso_11__9_, ADD_esteso_11__8_, ADD_esteso_11__7_,
         ADD_esteso_11__6_, ADD_esteso_11__5_, ADD_esteso_11__4_,
         ADD_esteso_11__3_, ADD_esteso_11__2_, ADD_esteso_11__1_,
         ADD_esteso_11__0_, ADD_esteso_12__17_, ADD_esteso_12__16_,
         ADD_esteso_12__15_, ADD_esteso_12__14_, ADD_esteso_12__13_,
         ADD_esteso_12__12_, ADD_esteso_12__11_, ADD_esteso_12__10_,
         ADD_esteso_12__9_, ADD_esteso_12__8_, ADD_esteso_12__7_,
         ADD_esteso_12__6_, ADD_esteso_12__5_, ADD_esteso_12__4_,
         ADD_esteso_12__3_, ADD_esteso_12__2_, ADD_esteso_12__1_,
         ADD_esteso_12__0_, ADD_esteso_13__17_, ADD_esteso_13__16_,
         ADD_esteso_13__15_, ADD_esteso_13__14_, ADD_esteso_13__13_,
         ADD_esteso_13__12_, ADD_esteso_13__11_, ADD_esteso_13__10_,
         ADD_esteso_13__9_, ADD_esteso_13__8_, ADD_esteso_13__7_,
         ADD_esteso_13__6_, ADD_esteso_13__5_, ADD_esteso_13__4_,
         ADD_esteso_13__3_, ADD_esteso_13__2_, ADD_esteso_13__1_,
         ADD_esteso_13__0_, ADD_esteso_14__17_, ADD_esteso_14__16_,
         ADD_esteso_14__15_, ADD_esteso_14__14_, ADD_esteso_14__13_,
         ADD_esteso_14__12_, ADD_esteso_14__11_, ADD_esteso_14__10_, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, ADD2_2_add_16_DP_OP_276_702_2_n50,
         ADD2_2_add_16_DP_OP_276_702_2_n49, ADD2_2_add_16_DP_OP_276_702_2_n48,
         ADD2_2_add_16_DP_OP_276_702_2_n47, ADD2_2_add_16_DP_OP_276_702_2_n46,
         ADD2_2_add_16_DP_OP_276_702_2_n45, ADD2_2_add_16_DP_OP_276_702_2_n44,
         ADD2_2_add_16_DP_OP_276_702_2_n43, ADD2_2_add_16_DP_OP_276_702_2_n42,
         ADD2_2_add_16_DP_OP_276_702_2_n41, ADD2_2_add_16_DP_OP_276_702_2_n40,
         ADD2_2_add_16_DP_OP_276_702_2_n39, ADD2_2_add_16_DP_OP_276_702_2_n38,
         ADD2_2_add_16_DP_OP_276_702_2_n37, ADD2_2_add_16_DP_OP_276_702_2_n36,
         ADD2_2_add_16_DP_OP_276_702_2_n35, ADD2_2_add_16_DP_OP_276_702_2_n34,
         ADD2_2_add_16_DP_OP_276_702_2_n33, ADD2_2_add_16_DP_OP_276_702_2_n32,
         ADD2_2_add_16_DP_OP_276_702_2_n31, ADD2_2_add_16_DP_OP_276_702_2_n30,
         ADD2_2_add_16_DP_OP_276_702_2_n29, ADD2_2_add_16_DP_OP_276_702_2_n28,
         ADD2_2_add_16_DP_OP_276_702_2_n27, ADD2_2_add_16_DP_OP_276_702_2_n26,
         ADD2_2_add_16_DP_OP_276_702_2_n25, ADD2_2_add_16_DP_OP_276_702_2_n24,
         ADD2_2_add_16_DP_OP_276_702_2_n23, ADD2_2_add_16_DP_OP_276_702_2_n22,
         ADD2_2_add_16_DP_OP_276_702_2_n21, ADD2_2_add_16_DP_OP_276_702_2_n20,
         ADD2_2_add_16_DP_OP_276_702_2_n19, ADD2_2_add_16_DP_OP_276_702_2_n18,
         ADD2_2_add_16_DP_OP_276_702_2_n17, ADD2_2_add_16_DP_OP_276_702_2_n16,
         ADD2_2_add_16_DP_OP_276_702_2_n15, ADD2_2_add_16_DP_OP_276_702_2_n14,
         ADD2_2_add_16_DP_OP_276_702_2_n13, ADD2_2_add_16_DP_OP_276_702_2_n12,
         ADD2_2_add_16_DP_OP_276_702_2_n11, ADD2_2_add_16_DP_OP_276_702_2_n10,
         ADD2_2_add_16_DP_OP_276_702_2_n9, ADD2_2_add_16_DP_OP_276_702_2_n8,
         ADD2_2_add_16_DP_OP_276_702_2_n7, ADD2_2_add_16_DP_OP_276_702_2_n6,
         ADD2_2_add_16_DP_OP_276_702_2_n5, ADD2_2_add_16_DP_OP_276_702_2_n4,
         ADD2_2_add_16_DP_OP_276_702_2_n3, ADD2_2_add_16_DP_OP_276_702_2_n2,
         ADD2_2_add_16_DP_OP_276_702_2_n1, ADD2_1_add_16_DP_OP_277_5600_1_n69,
         ADD2_1_add_16_DP_OP_277_5600_1_n68,
         ADD2_1_add_16_DP_OP_277_5600_1_n67,
         ADD2_1_add_16_DP_OP_277_5600_1_n66,
         ADD2_1_add_16_DP_OP_277_5600_1_n65,
         ADD2_1_add_16_DP_OP_277_5600_1_n64,
         ADD2_1_add_16_DP_OP_277_5600_1_n63,
         ADD2_1_add_16_DP_OP_277_5600_1_n62,
         ADD2_1_add_16_DP_OP_277_5600_1_n61,
         ADD2_1_add_16_DP_OP_277_5600_1_n60,
         ADD2_1_add_16_DP_OP_277_5600_1_n59,
         ADD2_1_add_16_DP_OP_277_5600_1_n58,
         ADD2_1_add_16_DP_OP_277_5600_1_n57,
         ADD2_1_add_16_DP_OP_277_5600_1_n56,
         ADD2_1_add_16_DP_OP_277_5600_1_n55,
         ADD2_1_add_16_DP_OP_277_5600_1_n54,
         ADD2_1_add_16_DP_OP_277_5600_1_n53,
         ADD2_1_add_16_DP_OP_277_5600_1_n52,
         ADD2_1_add_16_DP_OP_277_5600_1_n51,
         ADD2_1_add_16_DP_OP_277_5600_1_n50,
         ADD2_1_add_16_DP_OP_277_5600_1_n49,
         ADD2_1_add_16_DP_OP_277_5600_1_n48,
         ADD2_1_add_16_DP_OP_277_5600_1_n47,
         ADD2_1_add_16_DP_OP_277_5600_1_n46,
         ADD2_1_add_16_DP_OP_277_5600_1_n45,
         ADD2_1_add_16_DP_OP_277_5600_1_n44,
         ADD2_1_add_16_DP_OP_277_5600_1_n43,
         ADD2_1_add_16_DP_OP_277_5600_1_n42,
         ADD2_1_add_16_DP_OP_277_5600_1_n41,
         ADD2_1_add_16_DP_OP_277_5600_1_n40,
         ADD2_1_add_16_DP_OP_277_5600_1_n39,
         ADD2_1_add_16_DP_OP_277_5600_1_n38,
         ADD2_1_add_16_DP_OP_277_5600_1_n37,
         ADD2_1_add_16_DP_OP_277_5600_1_n36,
         ADD2_1_add_16_DP_OP_277_5600_1_n35,
         ADD2_1_add_16_DP_OP_277_5600_1_n34,
         ADD2_1_add_16_DP_OP_277_5600_1_n33,
         ADD2_1_add_16_DP_OP_277_5600_1_n32,
         ADD2_1_add_16_DP_OP_277_5600_1_n31,
         ADD2_1_add_16_DP_OP_277_5600_1_n30,
         ADD2_1_add_16_DP_OP_277_5600_1_n29,
         ADD2_1_add_16_DP_OP_277_5600_1_n28,
         ADD2_1_add_16_DP_OP_277_5600_1_n27,
         ADD2_1_add_16_DP_OP_277_5600_1_n26,
         ADD2_1_add_16_DP_OP_277_5600_1_n25,
         ADD2_1_add_16_DP_OP_277_5600_1_n24,
         ADD2_1_add_16_DP_OP_277_5600_1_n23,
         ADD2_1_add_16_DP_OP_277_5600_1_n22,
         ADD2_1_add_16_DP_OP_277_5600_1_n21,
         ADD2_1_add_16_DP_OP_277_5600_1_n20,
         ADD2_1_add_16_DP_OP_277_5600_1_n19,
         ADD2_1_add_16_DP_OP_277_5600_1_n18,
         ADD2_1_add_16_DP_OP_277_5600_1_n17,
         ADD2_1_add_16_DP_OP_277_5600_1_n16,
         ADD2_1_add_16_DP_OP_277_5600_1_n15,
         ADD2_1_add_16_DP_OP_277_5600_1_n14,
         ADD2_1_add_16_DP_OP_277_5600_1_n13,
         ADD2_1_add_16_DP_OP_277_5600_1_n12,
         ADD2_1_add_16_DP_OP_277_5600_1_n11,
         ADD2_1_add_16_DP_OP_277_5600_1_n10, ADD2_1_add_16_DP_OP_277_5600_1_n9,
         ADD2_1_add_16_DP_OP_277_5600_1_n8, ADD2_1_add_16_DP_OP_277_5600_1_n7,
         ADD2_1_add_16_DP_OP_277_5600_1_n6, ADD2_1_add_16_DP_OP_277_5600_1_n5,
         ADD2_1_add_16_DP_OP_277_5600_1_n4, ADD2_1_add_16_DP_OP_277_5600_1_n3,
         ADD2_1_add_16_DP_OP_277_5600_1_n2, ADD2_1_add_16_DP_OP_277_5600_1_n1,
         ADD3_1_add_16_carry_10_, ADD3_1_add_16_carry_11_,
         ADD3_1_add_16_carry_12_, ADD3_1_add_16_carry_13_,
         ADD3_1_add_16_carry_14_, ADD3_1_add_16_carry_15_,
         ADD3_1_add_16_carry_16_, ADD3_1_add_16_carry_17_, MULi_1_mult_15_n87,
         MULi_1_mult_15_n86, MULi_1_mult_15_n85, MULi_1_mult_15_n84,
         MULi_1_mult_15_n83, MULi_1_mult_15_n82, MULi_1_mult_15_n81,
         MULi_1_mult_15_n79, MULi_1_mult_15_n78, MULi_1_mult_15_n77,
         MULi_1_mult_15_n76, MULi_1_mult_15_n75, MULi_1_mult_15_n74,
         MULi_1_mult_15_n72, MULi_1_mult_15_n71, MULi_1_mult_15_n70,
         MULi_1_mult_15_n69, MULi_1_mult_15_n68, MULi_1_mult_15_n67,
         MULi_1_mult_15_n66, MULi_1_mult_15_n65, MULi_1_mult_15_n64,
         MULi_1_mult_15_n63, MULi_1_mult_15_n62, MULi_1_mult_15_n61,
         MULi_1_mult_15_n60, MULi_1_mult_15_n59, MULi_1_mult_15_n58,
         MULi_1_mult_15_n57, MULi_1_mult_15_n56, MULi_1_mult_15_n55,
         MULi_1_mult_15_n54, MULi_1_mult_15_n53, MULi_1_mult_15_n52,
         MULi_1_mult_15_n51, MULi_1_mult_15_n50, MULi_1_mult_15_n49,
         MULi_1_mult_15_n48, MULi_1_mult_15_n47, MULi_1_mult_15_n46,
         MULi_1_mult_15_n45, MULi_1_mult_15_n44, MULi_1_mult_15_n43,
         MULi_1_mult_15_n42, MULi_1_mult_15_n41, MULi_1_mult_15_n40,
         MULi_1_mult_15_n39, MULi_1_mult_15_n38, MULi_1_mult_15_n37,
         MULi_1_mult_15_n36, MULi_1_mult_15_n35, MULi_1_mult_15_n34,
         MULi_1_mult_15_n33, MULi_1_mult_15_n32, MULi_1_mult_15_n31,
         MULi_1_mult_15_n28, MULi_1_mult_15_n27, MULi_1_mult_15_n26,
         MULi_1_mult_15_n25, MULi_1_mult_15_n24, MULi_1_mult_15_n23,
         MULi_1_mult_15_n22, MULi_1_mult_15_n21, MULi_1_mult_15_n20,
         MULi_1_mult_15_n19, MULi_1_mult_15_n18, MULi_1_mult_15_n17,
         MULi_1_mult_15_n16, MULi_1_mult_15_n15, MULi_1_mult_15_n14,
         MULi_1_mult_15_n13, MULi_1_mult_15_n12, MULi_1_mult_15_n11,
         MULi_1_mult_15_n10, MULi_1_mult_15_n9, MULi_1_mult_15_n8,
         MULi_1_mult_15_n7, MULi_1_mult_15_n6, MULi_1_mult_15_n5,
         MULi_1_mult_15_n4, MULi_1_mult_15_n3, MULi_1_mult_15_n2,
         MULi_1_mult_15_n1, MULi_2_mult_15_n87, MULi_2_mult_15_n86,
         MULi_2_mult_15_n85, MULi_2_mult_15_n84, MULi_2_mult_15_n83,
         MULi_2_mult_15_n82, MULi_2_mult_15_n81, MULi_2_mult_15_n79,
         MULi_2_mult_15_n78, MULi_2_mult_15_n77, MULi_2_mult_15_n76,
         MULi_2_mult_15_n75, MULi_2_mult_15_n74, MULi_2_mult_15_n72,
         MULi_2_mult_15_n71, MULi_2_mult_15_n70, MULi_2_mult_15_n69,
         MULi_2_mult_15_n68, MULi_2_mult_15_n67, MULi_2_mult_15_n66,
         MULi_2_mult_15_n65, MULi_2_mult_15_n64, MULi_2_mult_15_n63,
         MULi_2_mult_15_n62, MULi_2_mult_15_n61, MULi_2_mult_15_n60,
         MULi_2_mult_15_n59, MULi_2_mult_15_n58, MULi_2_mult_15_n57,
         MULi_2_mult_15_n56, MULi_2_mult_15_n55, MULi_2_mult_15_n54,
         MULi_2_mult_15_n53, MULi_2_mult_15_n52, MULi_2_mult_15_n51,
         MULi_2_mult_15_n50, MULi_2_mult_15_n49, MULi_2_mult_15_n48,
         MULi_2_mult_15_n47, MULi_2_mult_15_n46, MULi_2_mult_15_n45,
         MULi_2_mult_15_n44, MULi_2_mult_15_n43, MULi_2_mult_15_n42,
         MULi_2_mult_15_n41, MULi_2_mult_15_n40, MULi_2_mult_15_n39,
         MULi_2_mult_15_n38, MULi_2_mult_15_n37, MULi_2_mult_15_n36,
         MULi_2_mult_15_n35, MULi_2_mult_15_n34, MULi_2_mult_15_n33,
         MULi_2_mult_15_n32, MULi_2_mult_15_n31, MULi_2_mult_15_n28,
         MULi_2_mult_15_n27, MULi_2_mult_15_n26, MULi_2_mult_15_n25,
         MULi_2_mult_15_n24, MULi_2_mult_15_n23, MULi_2_mult_15_n22,
         MULi_2_mult_15_n21, MULi_2_mult_15_n20, MULi_2_mult_15_n19,
         MULi_2_mult_15_n18, MULi_2_mult_15_n17, MULi_2_mult_15_n16,
         MULi_2_mult_15_n15, MULi_2_mult_15_n14, MULi_2_mult_15_n13,
         MULi_2_mult_15_n12, MULi_2_mult_15_n11, MULi_2_mult_15_n10,
         MULi_2_mult_15_n9, MULi_2_mult_15_n8, MULi_2_mult_15_n7,
         MULi_2_mult_15_n6, MULi_2_mult_15_n5, MULi_2_mult_15_n4,
         MULi_2_mult_15_n3, MULi_2_mult_15_n2, MULi_2_mult_15_n1,
         MULi_3_mult_15_n87, MULi_3_mult_15_n86, MULi_3_mult_15_n85,
         MULi_3_mult_15_n84, MULi_3_mult_15_n83, MULi_3_mult_15_n82,
         MULi_3_mult_15_n81, MULi_3_mult_15_n79, MULi_3_mult_15_n78,
         MULi_3_mult_15_n77, MULi_3_mult_15_n76, MULi_3_mult_15_n75,
         MULi_3_mult_15_n74, MULi_3_mult_15_n72, MULi_3_mult_15_n71,
         MULi_3_mult_15_n70, MULi_3_mult_15_n69, MULi_3_mult_15_n68,
         MULi_3_mult_15_n67, MULi_3_mult_15_n66, MULi_3_mult_15_n65,
         MULi_3_mult_15_n64, MULi_3_mult_15_n63, MULi_3_mult_15_n62,
         MULi_3_mult_15_n61, MULi_3_mult_15_n60, MULi_3_mult_15_n59,
         MULi_3_mult_15_n58, MULi_3_mult_15_n57, MULi_3_mult_15_n56,
         MULi_3_mult_15_n55, MULi_3_mult_15_n54, MULi_3_mult_15_n53,
         MULi_3_mult_15_n52, MULi_3_mult_15_n51, MULi_3_mult_15_n50,
         MULi_3_mult_15_n49, MULi_3_mult_15_n48, MULi_3_mult_15_n47,
         MULi_3_mult_15_n46, MULi_3_mult_15_n45, MULi_3_mult_15_n44,
         MULi_3_mult_15_n43, MULi_3_mult_15_n42, MULi_3_mult_15_n41,
         MULi_3_mult_15_n40, MULi_3_mult_15_n39, MULi_3_mult_15_n38,
         MULi_3_mult_15_n37, MULi_3_mult_15_n36, MULi_3_mult_15_n35,
         MULi_3_mult_15_n34, MULi_3_mult_15_n33, MULi_3_mult_15_n32,
         MULi_3_mult_15_n31, MULi_3_mult_15_n28, MULi_3_mult_15_n27,
         MULi_3_mult_15_n26, MULi_3_mult_15_n25, MULi_3_mult_15_n24,
         MULi_3_mult_15_n23, MULi_3_mult_15_n22, MULi_3_mult_15_n21,
         MULi_3_mult_15_n20, MULi_3_mult_15_n19, MULi_3_mult_15_n18,
         MULi_3_mult_15_n17, MULi_3_mult_15_n16, MULi_3_mult_15_n15,
         MULi_3_mult_15_n14, MULi_3_mult_15_n13, MULi_3_mult_15_n12,
         MULi_3_mult_15_n11, MULi_3_mult_15_n10, MULi_3_mult_15_n9,
         MULi_3_mult_15_n8, MULi_3_mult_15_n7, MULi_3_mult_15_n6,
         MULi_3_mult_15_n5, MULi_3_mult_15_n4, MULi_3_mult_15_n3,
         MULi_3_mult_15_n2, MULi_3_mult_15_n1, MULi_4_mult_15_n87,
         MULi_4_mult_15_n86, MULi_4_mult_15_n85, MULi_4_mult_15_n84,
         MULi_4_mult_15_n83, MULi_4_mult_15_n82, MULi_4_mult_15_n81,
         MULi_4_mult_15_n79, MULi_4_mult_15_n78, MULi_4_mult_15_n77,
         MULi_4_mult_15_n76, MULi_4_mult_15_n75, MULi_4_mult_15_n74,
         MULi_4_mult_15_n72, MULi_4_mult_15_n71, MULi_4_mult_15_n70,
         MULi_4_mult_15_n69, MULi_4_mult_15_n68, MULi_4_mult_15_n67,
         MULi_4_mult_15_n66, MULi_4_mult_15_n65, MULi_4_mult_15_n64,
         MULi_4_mult_15_n63, MULi_4_mult_15_n62, MULi_4_mult_15_n61,
         MULi_4_mult_15_n60, MULi_4_mult_15_n59, MULi_4_mult_15_n58,
         MULi_4_mult_15_n57, MULi_4_mult_15_n56, MULi_4_mult_15_n55,
         MULi_4_mult_15_n54, MULi_4_mult_15_n53, MULi_4_mult_15_n52,
         MULi_4_mult_15_n51, MULi_4_mult_15_n50, MULi_4_mult_15_n49,
         MULi_4_mult_15_n48, MULi_4_mult_15_n47, MULi_4_mult_15_n46,
         MULi_4_mult_15_n45, MULi_4_mult_15_n44, MULi_4_mult_15_n43,
         MULi_4_mult_15_n42, MULi_4_mult_15_n41, MULi_4_mult_15_n40,
         MULi_4_mult_15_n39, MULi_4_mult_15_n38, MULi_4_mult_15_n37,
         MULi_4_mult_15_n36, MULi_4_mult_15_n35, MULi_4_mult_15_n34,
         MULi_4_mult_15_n33, MULi_4_mult_15_n32, MULi_4_mult_15_n31,
         MULi_4_mult_15_n28, MULi_4_mult_15_n27, MULi_4_mult_15_n26,
         MULi_4_mult_15_n25, MULi_4_mult_15_n24, MULi_4_mult_15_n23,
         MULi_4_mult_15_n22, MULi_4_mult_15_n21, MULi_4_mult_15_n20,
         MULi_4_mult_15_n19, MULi_4_mult_15_n18, MULi_4_mult_15_n17,
         MULi_4_mult_15_n16, MULi_4_mult_15_n15, MULi_4_mult_15_n14,
         MULi_4_mult_15_n13, MULi_4_mult_15_n12, MULi_4_mult_15_n11,
         MULi_4_mult_15_n10, MULi_4_mult_15_n9, MULi_4_mult_15_n8,
         MULi_4_mult_15_n7, MULi_4_mult_15_n6, MULi_4_mult_15_n5,
         MULi_4_mult_15_n4, MULi_4_mult_15_n3, MULi_4_mult_15_n2,
         MULi_4_mult_15_n1, MULi_5_mult_15_n87, MULi_5_mult_15_n86,
         MULi_5_mult_15_n85, MULi_5_mult_15_n84, MULi_5_mult_15_n83,
         MULi_5_mult_15_n82, MULi_5_mult_15_n81, MULi_5_mult_15_n79,
         MULi_5_mult_15_n78, MULi_5_mult_15_n77, MULi_5_mult_15_n76,
         MULi_5_mult_15_n75, MULi_5_mult_15_n74, MULi_5_mult_15_n72,
         MULi_5_mult_15_n71, MULi_5_mult_15_n70, MULi_5_mult_15_n69,
         MULi_5_mult_15_n68, MULi_5_mult_15_n67, MULi_5_mult_15_n66,
         MULi_5_mult_15_n65, MULi_5_mult_15_n64, MULi_5_mult_15_n63,
         MULi_5_mult_15_n62, MULi_5_mult_15_n61, MULi_5_mult_15_n60,
         MULi_5_mult_15_n59, MULi_5_mult_15_n58, MULi_5_mult_15_n57,
         MULi_5_mult_15_n56, MULi_5_mult_15_n55, MULi_5_mult_15_n54,
         MULi_5_mult_15_n53, MULi_5_mult_15_n52, MULi_5_mult_15_n51,
         MULi_5_mult_15_n50, MULi_5_mult_15_n49, MULi_5_mult_15_n48,
         MULi_5_mult_15_n47, MULi_5_mult_15_n46, MULi_5_mult_15_n45,
         MULi_5_mult_15_n44, MULi_5_mult_15_n43, MULi_5_mult_15_n42,
         MULi_5_mult_15_n41, MULi_5_mult_15_n40, MULi_5_mult_15_n39,
         MULi_5_mult_15_n38, MULi_5_mult_15_n37, MULi_5_mult_15_n36,
         MULi_5_mult_15_n35, MULi_5_mult_15_n34, MULi_5_mult_15_n33,
         MULi_5_mult_15_n32, MULi_5_mult_15_n31, MULi_5_mult_15_n28,
         MULi_5_mult_15_n27, MULi_5_mult_15_n26, MULi_5_mult_15_n25,
         MULi_5_mult_15_n24, MULi_5_mult_15_n23, MULi_5_mult_15_n22,
         MULi_5_mult_15_n21, MULi_5_mult_15_n20, MULi_5_mult_15_n19,
         MULi_5_mult_15_n18, MULi_5_mult_15_n17, MULi_5_mult_15_n16,
         MULi_5_mult_15_n15, MULi_5_mult_15_n14, MULi_5_mult_15_n13,
         MULi_5_mult_15_n12, MULi_5_mult_15_n11, MULi_5_mult_15_n10,
         MULi_5_mult_15_n9, MULi_5_mult_15_n8, MULi_5_mult_15_n7,
         MULi_5_mult_15_n6, MULi_5_mult_15_n5, MULi_5_mult_15_n4,
         MULi_5_mult_15_n3, MULi_5_mult_15_n2, MULi_5_mult_15_n1,
         MULi_6_mult_15_n87, MULi_6_mult_15_n86, MULi_6_mult_15_n85,
         MULi_6_mult_15_n84, MULi_6_mult_15_n83, MULi_6_mult_15_n82,
         MULi_6_mult_15_n81, MULi_6_mult_15_n79, MULi_6_mult_15_n78,
         MULi_6_mult_15_n77, MULi_6_mult_15_n76, MULi_6_mult_15_n75,
         MULi_6_mult_15_n74, MULi_6_mult_15_n72, MULi_6_mult_15_n71,
         MULi_6_mult_15_n70, MULi_6_mult_15_n69, MULi_6_mult_15_n68,
         MULi_6_mult_15_n67, MULi_6_mult_15_n66, MULi_6_mult_15_n65,
         MULi_6_mult_15_n64, MULi_6_mult_15_n63, MULi_6_mult_15_n62,
         MULi_6_mult_15_n61, MULi_6_mult_15_n60, MULi_6_mult_15_n59,
         MULi_6_mult_15_n58, MULi_6_mult_15_n57, MULi_6_mult_15_n56,
         MULi_6_mult_15_n55, MULi_6_mult_15_n54, MULi_6_mult_15_n53,
         MULi_6_mult_15_n52, MULi_6_mult_15_n51, MULi_6_mult_15_n50,
         MULi_6_mult_15_n49, MULi_6_mult_15_n48, MULi_6_mult_15_n47,
         MULi_6_mult_15_n46, MULi_6_mult_15_n45, MULi_6_mult_15_n44,
         MULi_6_mult_15_n43, MULi_6_mult_15_n42, MULi_6_mult_15_n41,
         MULi_6_mult_15_n40, MULi_6_mult_15_n39, MULi_6_mult_15_n38,
         MULi_6_mult_15_n37, MULi_6_mult_15_n36, MULi_6_mult_15_n35,
         MULi_6_mult_15_n34, MULi_6_mult_15_n33, MULi_6_mult_15_n32,
         MULi_6_mult_15_n31, MULi_6_mult_15_n28, MULi_6_mult_15_n27,
         MULi_6_mult_15_n26, MULi_6_mult_15_n25, MULi_6_mult_15_n24,
         MULi_6_mult_15_n23, MULi_6_mult_15_n22, MULi_6_mult_15_n21,
         MULi_6_mult_15_n20, MULi_6_mult_15_n19, MULi_6_mult_15_n18,
         MULi_6_mult_15_n17, MULi_6_mult_15_n16, MULi_6_mult_15_n15,
         MULi_6_mult_15_n14, MULi_6_mult_15_n13, MULi_6_mult_15_n12,
         MULi_6_mult_15_n11, MULi_6_mult_15_n10, MULi_6_mult_15_n9,
         MULi_6_mult_15_n8, MULi_6_mult_15_n7, MULi_6_mult_15_n6,
         MULi_6_mult_15_n5, MULi_6_mult_15_n4, MULi_6_mult_15_n3,
         MULi_6_mult_15_n2, MULi_6_mult_15_n1, MULi_0_mult_15_n87,
         MULi_0_mult_15_n86, MULi_0_mult_15_n85, MULi_0_mult_15_n84,
         MULi_0_mult_15_n83, MULi_0_mult_15_n82, MULi_0_mult_15_n81,
         MULi_0_mult_15_n79, MULi_0_mult_15_n78, MULi_0_mult_15_n77,
         MULi_0_mult_15_n76, MULi_0_mult_15_n75, MULi_0_mult_15_n74,
         MULi_0_mult_15_n72, MULi_0_mult_15_n71, MULi_0_mult_15_n70,
         MULi_0_mult_15_n69, MULi_0_mult_15_n68, MULi_0_mult_15_n67,
         MULi_0_mult_15_n66, MULi_0_mult_15_n65, MULi_0_mult_15_n64,
         MULi_0_mult_15_n63, MULi_0_mult_15_n62, MULi_0_mult_15_n61,
         MULi_0_mult_15_n60, MULi_0_mult_15_n59, MULi_0_mult_15_n58,
         MULi_0_mult_15_n57, MULi_0_mult_15_n56, MULi_0_mult_15_n55,
         MULi_0_mult_15_n54, MULi_0_mult_15_n53, MULi_0_mult_15_n52,
         MULi_0_mult_15_n51, MULi_0_mult_15_n50, MULi_0_mult_15_n49,
         MULi_0_mult_15_n48, MULi_0_mult_15_n47, MULi_0_mult_15_n46,
         MULi_0_mult_15_n45, MULi_0_mult_15_n44, MULi_0_mult_15_n43,
         MULi_0_mult_15_n42, MULi_0_mult_15_n41, MULi_0_mult_15_n40,
         MULi_0_mult_15_n39, MULi_0_mult_15_n38, MULi_0_mult_15_n37,
         MULi_0_mult_15_n36, MULi_0_mult_15_n35, MULi_0_mult_15_n34,
         MULi_0_mult_15_n33, MULi_0_mult_15_n32, MULi_0_mult_15_n31,
         MULi_0_mult_15_n28, MULi_0_mult_15_n27, MULi_0_mult_15_n26,
         MULi_0_mult_15_n25, MULi_0_mult_15_n24, MULi_0_mult_15_n23,
         MULi_0_mult_15_n22, MULi_0_mult_15_n21, MULi_0_mult_15_n20,
         MULi_0_mult_15_n19, MULi_0_mult_15_n18, MULi_0_mult_15_n17,
         MULi_0_mult_15_n16, MULi_0_mult_15_n15, MULi_0_mult_15_n14,
         MULi_0_mult_15_n13, MULi_0_mult_15_n12, MULi_0_mult_15_n11,
         MULi_0_mult_15_n10, MULi_0_mult_15_n9, MULi_0_mult_15_n8,
         MULi_0_mult_15_n7, MULi_0_mult_15_n6, MULi_0_mult_15_n5,
         MULi_0_mult_15_n4, MULi_0_mult_15_n3, MULi_0_mult_15_n2,
         MULi_0_mult_15_n1, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690;
  wire   [55:0] SR_to_MUL;
  wire   [55:0] TEMP_H;
  wire   [111:0] MUL_to_PIPE1;
  wire   [5:0] SR_SRI_bit_temp_out;

  DFFRQX2 REG_OUT_VIN_q_reg ( .D(PIPE2_to_REGOUT), .CK(CLK), .RN(RST_n), .Q(
        VOUT) );
  DFFRQX2 REG_OUT_q_reg_0_ ( .D(ADD_esteso_14__10_), .CK(CLK), .RN(RST_n), .Q(
        DOUT[0]) );
  DFFRQX2 REG_OUT_q_reg_1_ ( .D(ADD_esteso_14__11_), .CK(CLK), .RN(RST_n), .Q(
        DOUT[1]) );
  DFFRQX2 REG_OUT_q_reg_2_ ( .D(ADD_esteso_14__12_), .CK(CLK), .RN(RST_n), .Q(
        DOUT[2]) );
  DFFRQX2 REG_OUT_q_reg_3_ ( .D(ADD_esteso_14__13_), .CK(CLK), .RN(RST_n), .Q(
        DOUT[3]) );
  DFFRQX2 REG_OUT_q_reg_4_ ( .D(ADD_esteso_14__14_), .CK(CLK), .RN(RST_n), .Q(
        DOUT[4]) );
  DFFRQX2 REG_OUT_q_reg_5_ ( .D(ADD_esteso_14__15_), .CK(CLK), .RN(RST_n), .Q(
        DOUT[5]) );
  DFFRQX2 REG_OUT_q_reg_6_ ( .D(ADD_esteso_14__16_), .CK(CLK), .RN(RST_n), .Q(
        DOUT[6]) );
  DFFRQX2 REG_OUT_q_reg_7_ ( .D(ADD_esteso_14__17_), .CK(CLK), .RN(RST_n), .Q(
        DOUT[7]) );
  DFFRQX2 PIPE1_VIN_q_reg ( .D(MUX_to_PIPE1), .CK(CLK), .RN(RST_n), .Q(
        PIPE1_to_PIPE2) );
  DFFRQX2 PIPE2_VIN_q_reg ( .D(PIPE1_to_PIPE2), .CK(CLK), .RN(RST_n), .Q(
        PIPE2_to_REGOUT) );
  DFFRQX2 PIPE2_1_q_reg_10_ ( .D(ADD_esteso_10__10_), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_12__10_) );
  DFFRQX2 PIPE2_1_q_reg_11_ ( .D(ADD_esteso_10__11_), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_12__11_) );
  DFFRQX2 PIPE2_1_q_reg_12_ ( .D(ADD_esteso_10__12_), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_12__12_) );
  DFFRQX2 PIPE2_1_q_reg_13_ ( .D(ADD_esteso_10__13_), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_12__13_) );
  DFFRQX2 PIPE2_1_q_reg_14_ ( .D(ADD_esteso_10__14_), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_12__14_) );
  DFFRQX2 PIPE2_1_q_reg_15_ ( .D(ADD_esteso_10__15_), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_12__15_) );
  DFFRQX2 PIPE2_1_q_reg_16_ ( .D(ADD_esteso_10__16_), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_12__16_) );
  DFFRQX2 PIPE2_1_q_reg_17_ ( .D(ADD_esteso_10__17_), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_12__17_) );
  DFFRQX2 PIPE2_2_q_reg_10_ ( .D(ADD_esteso_11__10_), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_13__10_) );
  DFFRQX2 PIPE2_2_q_reg_11_ ( .D(ADD_esteso_11__11_), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_13__11_) );
  DFFRQX2 PIPE2_2_q_reg_12_ ( .D(ADD_esteso_11__12_), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_13__12_) );
  DFFRQX2 PIPE2_2_q_reg_13_ ( .D(ADD_esteso_11__13_), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_13__13_) );
  DFFRQX2 PIPE2_2_q_reg_14_ ( .D(ADD_esteso_11__14_), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_13__14_) );
  DFFRQX2 PIPE2_2_q_reg_15_ ( .D(ADD_esteso_11__15_), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_13__15_) );
  DFFRQX2 PIPE2_2_q_reg_16_ ( .D(ADD_esteso_11__16_), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_13__16_) );
  DFFRQX2 PIPE2_2_q_reg_17_ ( .D(ADD_esteso_11__17_), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_13__17_) );
  DFFRQX2 SR_SRI_bit_regi_0_q_reg ( .D(n61), .CK(CLK), .RN(RST_n), .Q(
        SR_SRI_bit_temp_out[1]) );
  DFFRQX2 SR_SRI_bit_regi_1_q_reg ( .D(n60), .CK(CLK), .RN(RST_n), .Q(
        SR_SRI_bit_temp_out[2]) );
  DFFRQX2 SR_SRI_bit_regi_2_q_reg ( .D(n59), .CK(CLK), .RN(RST_n), .Q(
        SR_SRI_bit_temp_out[3]) );
  DFFRQX2 SR_SRI_bit_regi_3_q_reg ( .D(n58), .CK(CLK), .RN(RST_n), .Q(
        SR_SRI_bit_temp_out[4]) );
  DFFRQX2 SR_SRI_bit_regi_4_q_reg ( .D(n57), .CK(CLK), .RN(RST_n), .Q(
        SR_SRI_bit_temp_out[5]) );
  DFFRQX2 PIPE1_i_5_q_reg_15_ ( .D(MUL_to_PIPE1[31]), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_5__17_) );
  DFFRQX2 SR_SRI_bit_regi_5_q_reg ( .D(n56), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUX) );
  DFFRQX2 SR_SRI_bit_reg0_q_reg ( .D(n62), .CK(CLK), .RN(RST_n), .Q(
        SR_SRI_bit_temp_out[0]) );
  DFFRQX2 PIPE1_i_0_q_reg_15_ ( .D(MUL_to_PIPE1[111]), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_0__17_) );
  DFFRQX2 PIPE1_i_6_q_reg_15_ ( .D(MUL_to_PIPE1[15]), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_6__17_) );
  DFFRQX2 PIPE1_i_4_q_reg_15_ ( .D(MUL_to_PIPE1[47]), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_4__17_) );
  DFFRQX2 PIPE1_i_3_q_reg_15_ ( .D(MUL_to_PIPE1[63]), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_3__17_) );
  DFFRQX2 PIPE1_i_2_q_reg_15_ ( .D(MUL_to_PIPE1[79]), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_2__17_) );
  DFFRQX2 PIPE1_i_1_q_reg_15_ ( .D(MUL_to_PIPE1[95]), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_1__17_) );
  DFFRQX2 PIPE1_i_6_q_reg_10_ ( .D(MUL_to_PIPE1[10]), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_6__10_) );
  DFFRQX2 PIPE1_i_6_q_reg_11_ ( .D(MUL_to_PIPE1[11]), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_6__11_) );
  DFFRQX2 PIPE1_i_6_q_reg_12_ ( .D(MUL_to_PIPE1[12]), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_6__12_) );
  DFFRQX2 PIPE1_i_6_q_reg_13_ ( .D(MUL_to_PIPE1[13]), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_6__13_) );
  DFFRQX2 PIPE1_i_6_q_reg_14_ ( .D(MUL_to_PIPE1[14]), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_6__14_) );
  DFFRQX2 PIPE1_i_5_q_reg_10_ ( .D(MUL_to_PIPE1[26]), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_5__10_) );
  DFFRQX2 PIPE1_i_5_q_reg_11_ ( .D(MUL_to_PIPE1[27]), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_5__11_) );
  DFFRQX2 PIPE1_i_5_q_reg_12_ ( .D(MUL_to_PIPE1[28]), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_5__12_) );
  DFFRQX2 PIPE1_i_5_q_reg_13_ ( .D(MUL_to_PIPE1[29]), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_5__13_) );
  DFFRQX2 PIPE1_i_5_q_reg_14_ ( .D(MUL_to_PIPE1[30]), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_5__14_) );
  DFFRQX2 PIPE1_i_4_q_reg_10_ ( .D(MUL_to_PIPE1[42]), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_4__10_) );
  DFFRQX2 PIPE1_i_4_q_reg_11_ ( .D(MUL_to_PIPE1[43]), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_4__11_) );
  DFFRQX2 PIPE1_i_4_q_reg_12_ ( .D(MUL_to_PIPE1[44]), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_4__12_) );
  DFFRQX2 PIPE1_i_4_q_reg_13_ ( .D(MUL_to_PIPE1[45]), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_4__13_) );
  DFFRQX2 PIPE1_i_4_q_reg_14_ ( .D(MUL_to_PIPE1[46]), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_4__14_) );
  DFFRQX2 PIPE1_i_2_q_reg_10_ ( .D(MUL_to_PIPE1[74]), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_2__10_) );
  DFFRQX2 PIPE1_i_2_q_reg_11_ ( .D(MUL_to_PIPE1[75]), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_2__11_) );
  DFFRQX2 PIPE1_i_2_q_reg_12_ ( .D(MUL_to_PIPE1[76]), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_2__12_) );
  DFFRQX2 PIPE1_i_2_q_reg_13_ ( .D(MUL_to_PIPE1[77]), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_2__13_) );
  DFFRQX2 PIPE1_i_2_q_reg_14_ ( .D(MUL_to_PIPE1[78]), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_2__14_) );
  DFFRQX2 PIPE1_i_0_q_reg_10_ ( .D(MUL_to_PIPE1[106]), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_0__10_) );
  DFFRQX2 PIPE1_i_0_q_reg_11_ ( .D(MUL_to_PIPE1[107]), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_0__11_) );
  DFFRQX2 PIPE1_i_0_q_reg_12_ ( .D(MUL_to_PIPE1[108]), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_0__12_) );
  DFFRQX2 PIPE1_i_0_q_reg_13_ ( .D(MUL_to_PIPE1[109]), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_0__13_) );
  DFFRQX2 PIPE1_i_0_q_reg_14_ ( .D(MUL_to_PIPE1[110]), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_0__14_) );
  DFFRQX2 PIPE1_i_1_q_reg_10_ ( .D(MUL_to_PIPE1[90]), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_1__10_) );
  DFFRQX2 PIPE1_i_1_q_reg_11_ ( .D(MUL_to_PIPE1[91]), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_1__11_) );
  DFFRQX2 PIPE1_i_1_q_reg_12_ ( .D(MUL_to_PIPE1[92]), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_1__12_) );
  DFFRQX2 PIPE1_i_1_q_reg_13_ ( .D(MUL_to_PIPE1[93]), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_1__13_) );
  DFFRQX2 PIPE1_i_1_q_reg_14_ ( .D(MUL_to_PIPE1[94]), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_1__14_) );
  DFFRQX2 PIPE1_i_3_q_reg_10_ ( .D(MUL_to_PIPE1[58]), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_3__10_) );
  DFFRQX2 PIPE1_i_3_q_reg_11_ ( .D(MUL_to_PIPE1[59]), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_3__11_) );
  DFFRQX2 PIPE1_i_3_q_reg_12_ ( .D(MUL_to_PIPE1[60]), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_3__12_) );
  DFFRQX2 PIPE1_i_3_q_reg_13_ ( .D(MUL_to_PIPE1[61]), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_3__13_) );
  DFFRQX2 PIPE1_i_3_q_reg_14_ ( .D(MUL_to_PIPE1[62]), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_3__14_) );
  DFFRQX2 PIPE2_2_q_reg_8_ ( .D(ADD_esteso_11__8_), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_13__8_) );
  DFFRQX2 PIPE2_1_q_reg_9_ ( .D(ADD_esteso_10__9_), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_12__9_) );
  DFFRQX2 PIPE2_1_q_reg_8_ ( .D(ADD_esteso_10__8_), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_12__8_) );
  DFFRQX2 PIPE2_2_q_reg_9_ ( .D(ADD_esteso_11__9_), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_13__9_) );
  DFFRQX2 PIPE1_i_6_q_reg_5_ ( .D(MUL_to_PIPE1[5]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_6__5_) );
  DFFRQX2 PIPE1_i_6_q_reg_6_ ( .D(MUL_to_PIPE1[6]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_6__6_) );
  DFFRQX2 PIPE1_i_6_q_reg_7_ ( .D(MUL_to_PIPE1[7]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_6__7_) );
  DFFRQX2 PIPE1_i_6_q_reg_8_ ( .D(MUL_to_PIPE1[8]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_6__8_) );
  DFFRQX2 PIPE1_i_6_q_reg_9_ ( .D(MUL_to_PIPE1[9]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_6__9_) );
  DFFRQX2 PIPE1_i_5_q_reg_5_ ( .D(MUL_to_PIPE1[21]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_5__5_) );
  DFFRQX2 PIPE1_i_5_q_reg_6_ ( .D(MUL_to_PIPE1[22]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_5__6_) );
  DFFRQX2 PIPE1_i_5_q_reg_7_ ( .D(MUL_to_PIPE1[23]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_5__7_) );
  DFFRQX2 PIPE1_i_5_q_reg_8_ ( .D(MUL_to_PIPE1[24]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_5__8_) );
  DFFRQX2 PIPE1_i_5_q_reg_9_ ( .D(MUL_to_PIPE1[25]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_5__9_) );
  DFFRQX2 PIPE1_i_4_q_reg_4_ ( .D(MUL_to_PIPE1[36]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_4__4_) );
  DFFRQX2 PIPE1_i_4_q_reg_5_ ( .D(MUL_to_PIPE1[37]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_4__5_) );
  DFFRQX2 PIPE1_i_4_q_reg_6_ ( .D(MUL_to_PIPE1[38]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_4__6_) );
  DFFRQX2 PIPE1_i_4_q_reg_7_ ( .D(MUL_to_PIPE1[39]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_4__7_) );
  DFFRQX2 PIPE1_i_4_q_reg_8_ ( .D(MUL_to_PIPE1[40]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_4__8_) );
  DFFRQX2 PIPE1_i_4_q_reg_9_ ( .D(MUL_to_PIPE1[41]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_4__9_) );
  DFFRQX2 PIPE1_i_2_q_reg_5_ ( .D(MUL_to_PIPE1[69]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_2__5_) );
  DFFRQX2 PIPE1_i_2_q_reg_6_ ( .D(MUL_to_PIPE1[70]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_2__6_) );
  DFFRQX2 PIPE1_i_2_q_reg_7_ ( .D(MUL_to_PIPE1[71]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_2__7_) );
  DFFRQX2 PIPE1_i_2_q_reg_8_ ( .D(MUL_to_PIPE1[72]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_2__8_) );
  DFFRQX2 PIPE1_i_2_q_reg_9_ ( .D(MUL_to_PIPE1[73]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_2__9_) );
  DFFRQX2 PIPE1_i_0_q_reg_5_ ( .D(MUL_to_PIPE1[101]), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_0__5_) );
  DFFRQX2 PIPE1_i_0_q_reg_6_ ( .D(MUL_to_PIPE1[102]), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_0__6_) );
  DFFRQX2 PIPE1_i_0_q_reg_7_ ( .D(MUL_to_PIPE1[103]), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_0__7_) );
  DFFRQX2 PIPE1_i_0_q_reg_8_ ( .D(MUL_to_PIPE1[104]), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_0__8_) );
  DFFRQX2 PIPE1_i_0_q_reg_9_ ( .D(MUL_to_PIPE1[105]), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_0__9_) );
  DFFRQX2 PIPE1_i_1_q_reg_5_ ( .D(MUL_to_PIPE1[85]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_1__5_) );
  DFFRQX2 PIPE1_i_1_q_reg_6_ ( .D(MUL_to_PIPE1[86]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_1__6_) );
  DFFRQX2 PIPE1_i_1_q_reg_7_ ( .D(MUL_to_PIPE1[87]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_1__7_) );
  DFFRQX2 PIPE1_i_1_q_reg_8_ ( .D(MUL_to_PIPE1[88]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_1__8_) );
  DFFRQX2 PIPE1_i_1_q_reg_9_ ( .D(MUL_to_PIPE1[89]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_1__9_) );
  DFFRQX2 PIPE1_i_3_q_reg_5_ ( .D(MUL_to_PIPE1[53]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_3__5_) );
  DFFRQX2 PIPE1_i_3_q_reg_6_ ( .D(MUL_to_PIPE1[54]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_3__6_) );
  DFFRQX2 PIPE1_i_3_q_reg_7_ ( .D(MUL_to_PIPE1[55]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_3__7_) );
  DFFRQX2 PIPE1_i_3_q_reg_8_ ( .D(MUL_to_PIPE1[56]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_3__8_) );
  DFFRQX2 PIPE1_i_3_q_reg_9_ ( .D(MUL_to_PIPE1[57]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_3__9_) );
  DFFRQX2 PIPE2_2_q_reg_6_ ( .D(ADD_esteso_11__6_), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_13__6_) );
  DFFRQX2 PIPE2_1_q_reg_5_ ( .D(ADD_esteso_10__5_), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_12__5_) );
  DFFRQX2 PIPE2_1_q_reg_7_ ( .D(ADD_esteso_10__7_), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_12__7_) );
  DFFRQX2 PIPE2_1_q_reg_6_ ( .D(ADD_esteso_10__6_), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_12__6_) );
  DFFRQX2 PIPE2_2_q_reg_5_ ( .D(ADD_esteso_11__5_), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_13__5_) );
  DFFRQX2 PIPE2_2_q_reg_7_ ( .D(ADD_esteso_11__7_), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_13__7_) );
  DFFRQX2 SR_SRI_regi_6_q_reg_7_ ( .D(n8), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[7]) );
  DFFRQX2 PIPE1_i_4_q_reg_1_ ( .D(MUL_to_PIPE1[33]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_4__1_) );
  DFFRQX2 PIPE1_i_3_q_reg_1_ ( .D(MUL_to_PIPE1[49]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_3__1_) );
  DFFRQX2 PIPE1_i_2_q_reg_0_ ( .D(MUL_to_PIPE1[64]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_2__0_) );
  DFFRQX2 PIPE1_i_0_q_reg_1_ ( .D(MUL_to_PIPE1[97]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_0__1_) );
  DFFRQX2 PIPE1_i_6_q_reg_2_ ( .D(MUL_to_PIPE1[2]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_6__2_) );
  DFFRQX2 PIPE1_i_6_q_reg_3_ ( .D(MUL_to_PIPE1[3]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_6__3_) );
  DFFRQX2 PIPE1_i_6_q_reg_4_ ( .D(MUL_to_PIPE1[4]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_6__4_) );
  DFFRQX2 PIPE1_i_5_q_reg_0_ ( .D(MUL_to_PIPE1[16]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_5__0_) );
  DFFRQX2 PIPE1_i_3_q_reg_0_ ( .D(MUL_to_PIPE1[48]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_3__0_) );
  DFFRQX2 PIPE1_i_0_q_reg_0_ ( .D(MUL_to_PIPE1[96]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_0__0_) );
  DFFRQX2 PIPE1_i_6_q_reg_1_ ( .D(MUL_to_PIPE1[1]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_6__1_) );
  DFFRQX2 PIPE1_i_5_q_reg_2_ ( .D(MUL_to_PIPE1[18]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_5__2_) );
  DFFRQX2 PIPE1_i_5_q_reg_3_ ( .D(MUL_to_PIPE1[19]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_5__3_) );
  DFFRQX2 PIPE1_i_5_q_reg_4_ ( .D(MUL_to_PIPE1[20]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_5__4_) );
  DFFRQX2 PIPE1_i_4_q_reg_0_ ( .D(MUL_to_PIPE1[32]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_4__0_) );
  DFFRQX2 PIPE1_i_2_q_reg_1_ ( .D(MUL_to_PIPE1[65]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_2__1_) );
  DFFRQX2 PIPE1_i_6_q_reg_0_ ( .D(MUL_to_PIPE1[0]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_6__0_) );
  DFFRQX2 PIPE1_i_4_q_reg_2_ ( .D(MUL_to_PIPE1[34]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_4__2_) );
  DFFRQX2 PIPE1_i_4_q_reg_3_ ( .D(MUL_to_PIPE1[35]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_4__3_) );
  DFFRQX2 PIPE1_i_2_q_reg_2_ ( .D(MUL_to_PIPE1[66]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_2__2_) );
  DFFRQX2 PIPE1_i_2_q_reg_3_ ( .D(MUL_to_PIPE1[67]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_2__3_) );
  DFFRQX2 PIPE1_i_2_q_reg_4_ ( .D(MUL_to_PIPE1[68]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_2__4_) );
  DFFRQX2 PIPE1_i_5_q_reg_1_ ( .D(MUL_to_PIPE1[17]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_5__1_) );
  DFFRQX2 PIPE1_i_1_q_reg_0_ ( .D(MUL_to_PIPE1[80]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_1__0_) );
  DFFRQX2 PIPE1_i_1_q_reg_1_ ( .D(MUL_to_PIPE1[81]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_1__1_) );
  DFFRQX2 PIPE1_i_0_q_reg_2_ ( .D(MUL_to_PIPE1[98]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_0__2_) );
  DFFRQX2 PIPE1_i_0_q_reg_3_ ( .D(MUL_to_PIPE1[99]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_0__3_) );
  DFFRQX2 PIPE1_i_0_q_reg_4_ ( .D(MUL_to_PIPE1[100]), .CK(CLK), .RN(RST_n), 
        .Q(ADD_esteso_0__4_) );
  DFFRQX2 PIPE1_i_1_q_reg_2_ ( .D(MUL_to_PIPE1[82]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_1__2_) );
  DFFRQX2 PIPE1_i_1_q_reg_3_ ( .D(MUL_to_PIPE1[83]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_1__3_) );
  DFFRQX2 PIPE1_i_1_q_reg_4_ ( .D(MUL_to_PIPE1[84]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_1__4_) );
  DFFRQX2 PIPE1_i_3_q_reg_2_ ( .D(MUL_to_PIPE1[50]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_3__2_) );
  DFFRQX2 PIPE1_i_3_q_reg_3_ ( .D(MUL_to_PIPE1[51]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_3__3_) );
  DFFRQX2 PIPE1_i_3_q_reg_4_ ( .D(MUL_to_PIPE1[52]), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_3__4_) );
  DFFRQX2 PIPE2_2_q_reg_2_ ( .D(ADD_esteso_11__2_), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_13__2_) );
  DFFRQX2 PIPE2_2_q_reg_4_ ( .D(ADD_esteso_11__4_), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_13__4_) );
  DFFRQX2 PIPE2_1_q_reg_3_ ( .D(ADD_esteso_10__3_), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_12__3_) );
  DFFRQX2 PIPE2_1_q_reg_2_ ( .D(ADD_esteso_10__2_), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_12__2_) );
  DFFRQX2 PIPE2_1_q_reg_4_ ( .D(ADD_esteso_10__4_), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_12__4_) );
  DFFRQX2 PIPE2_2_q_reg_3_ ( .D(ADD_esteso_11__3_), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_13__3_) );
  DFFRQX2 SR_SRI_regi_6_q_reg_5_ ( .D(n20), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[5]) );
  DFFRQX2 PIPE2_1_q_reg_0_ ( .D(ADD_esteso_10__0_), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_12__0_) );
  DFFRQX2 PIPE2_2_q_reg_0_ ( .D(ADD_esteso_11__0_), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_13__0_) );
  DFFRQX2 PIPE2_2_q_reg_1_ ( .D(ADD_esteso_11__1_), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_13__1_) );
  DFFRQX2 PIPE2_1_q_reg_1_ ( .D(ADD_esteso_10__1_), .CK(CLK), .RN(RST_n), .Q(
        ADD_esteso_12__1_) );
  DFFRQX2 SR_SRI_regi_6_q_reg_3_ ( .D(n32), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[3]) );
  DFFRQX2 SR_SRI_regi_6_q_reg_1_ ( .D(n44), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[1]) );
  MX2X1 U50 ( .A(n114), .B(n116), .S0(VIN), .Y(n55) );
  MX2X1 U46 ( .A(n115), .B(n113), .S0(VIN), .Y(n51) );
  MX2X1 U48 ( .A(n111), .B(n112), .S0(VIN), .Y(n53) );
  MX2X1 U49 ( .A(n112), .B(n114), .S0(VIN), .Y(n54) );
  MX2X1 U45 ( .A(n103), .B(n115), .S0(VIN), .Y(n50) );
  MX2X1 U47 ( .A(n113), .B(n111), .S0(VIN), .Y(n52) );
  MX2X1 U65 ( .A(n116), .B(DIN[0]), .S0(VIN), .Y(n70) );
  MX2X1 U33 ( .A(SR_to_MUL[2]), .B(SR_to_MUL[10]), .S0(VIN), .Y(n38) );
  MX2X1 U35 ( .A(SR_to_MUL[18]), .B(SR_to_MUL[26]), .S0(VIN), .Y(n40) );
  MX2X1 U37 ( .A(SR_to_MUL[34]), .B(SR_to_MUL[42]), .S0(VIN), .Y(n42) );
  MX2X1 U34 ( .A(SR_to_MUL[10]), .B(SR_to_MUL[18]), .S0(VIN), .Y(n39) );
  MX2X1 U38 ( .A(SR_to_MUL[42]), .B(SR_to_MUL[50]), .S0(VIN), .Y(n43) );
  MX2X1 U36 ( .A(SR_to_MUL[26]), .B(SR_to_MUL[34]), .S0(VIN), .Y(n41) );
  MX2X1 U12 ( .A(SR_to_MUL[30]), .B(SR_to_MUL[38]), .S0(VIN), .Y(n17) );
  MX2X1 U25 ( .A(SR_to_MUL[36]), .B(SR_to_MUL[44]), .S0(VIN), .Y(n30) );
  MX2X1 U26 ( .A(SR_to_MUL[44]), .B(SR_to_MUL[52]), .S0(VIN), .Y(n31) );
  MX2X1 U23 ( .A(SR_to_MUL[20]), .B(SR_to_MUL[28]), .S0(VIN), .Y(n28) );
  MX2X1 U21 ( .A(SR_to_MUL[4]), .B(SR_to_MUL[12]), .S0(VIN), .Y(n26) );
  MX2X1 U9 ( .A(SR_to_MUL[6]), .B(SR_to_MUL[14]), .S0(VIN), .Y(n14) );
  MX2X1 U11 ( .A(SR_to_MUL[22]), .B(SR_to_MUL[30]), .S0(VIN), .Y(n16) );
  MX2X1 U24 ( .A(SR_to_MUL[28]), .B(SR_to_MUL[36]), .S0(VIN), .Y(n29) );
  MX2X1 U13 ( .A(SR_to_MUL[38]), .B(SR_to_MUL[46]), .S0(VIN), .Y(n18) );
  MX2X1 U22 ( .A(SR_to_MUL[12]), .B(SR_to_MUL[20]), .S0(VIN), .Y(n27) );
  MX2X1 U14 ( .A(SR_to_MUL[46]), .B(SR_to_MUL[54]), .S0(VIN), .Y(n19) );
  MX2X1 U10 ( .A(SR_to_MUL[14]), .B(SR_to_MUL[22]), .S0(VIN), .Y(n15) );
  MX2X1 U61 ( .A(SR_to_MUL[52]), .B(DIN[4]), .S0(VIN), .Y(n66) );
  MX2X1 U59 ( .A(SR_to_MUL[54]), .B(DIN[6]), .S0(VIN), .Y(n64) );
  MX2X1 U63 ( .A(SR_to_MUL[50]), .B(DIN[2]), .S0(VIN), .Y(n68) );
  MX2X1 U64 ( .A(SR_to_MUL[49]), .B(DIN[1]), .S0(VIN), .Y(n69) );
  MX2X1 U62 ( .A(SR_to_MUL[51]), .B(DIN[3]), .S0(VIN), .Y(n67) );
  MX2X1 U60 ( .A(SR_to_MUL[53]), .B(DIN[5]), .S0(VIN), .Y(n65) );
  MX2X1 U58 ( .A(SR_to_MUL[55]), .B(DIN[7]), .S0(VIN), .Y(n63) );
  MX2X1 U2 ( .A(SR_to_MUL[7]), .B(SR_to_MUL[15]), .S0(VIN), .Y(n8) );
  MX2X1 U31 ( .A(SR_to_MUL[35]), .B(SR_to_MUL[43]), .S0(VIN), .Y(n36) );
  MX2X1 U42 ( .A(SR_to_MUL[25]), .B(SR_to_MUL[33]), .S0(VIN), .Y(n47) );
  MX2X1 U17 ( .A(SR_to_MUL[21]), .B(SR_to_MUL[29]), .S0(VIN), .Y(n22) );
  MX2X1 U43 ( .A(SR_to_MUL[33]), .B(SR_to_MUL[41]), .S0(VIN), .Y(n48) );
  MX2X1 U19 ( .A(SR_to_MUL[37]), .B(SR_to_MUL[45]), .S0(VIN), .Y(n24) );
  MX2X1 U20 ( .A(SR_to_MUL[45]), .B(SR_to_MUL[53]), .S0(VIN), .Y(n25) );
  MX2X1 U41 ( .A(SR_to_MUL[17]), .B(SR_to_MUL[25]), .S0(VIN), .Y(n46) );
  MX2X1 U40 ( .A(SR_to_MUL[9]), .B(SR_to_MUL[17]), .S0(VIN), .Y(n45) );
  MX2X1 U27 ( .A(SR_to_MUL[3]), .B(SR_to_MUL[11]), .S0(VIN), .Y(n32) );
  MX2X1 U29 ( .A(SR_to_MUL[19]), .B(SR_to_MUL[27]), .S0(VIN), .Y(n34) );
  MX2X1 U30 ( .A(SR_to_MUL[27]), .B(SR_to_MUL[35]), .S0(VIN), .Y(n35) );
  MX2X1 U28 ( .A(SR_to_MUL[11]), .B(SR_to_MUL[19]), .S0(VIN), .Y(n33) );
  MX2X1 U39 ( .A(SR_to_MUL[1]), .B(SR_to_MUL[9]), .S0(VIN), .Y(n44) );
  MX2X1 U5 ( .A(SR_to_MUL[23]), .B(SR_to_MUL[31]), .S0(VIN), .Y(n10) );
  MX2X1 U16 ( .A(SR_to_MUL[13]), .B(SR_to_MUL[21]), .S0(VIN), .Y(n21) );
  MX2X1 U32 ( .A(SR_to_MUL[43]), .B(SR_to_MUL[51]), .S0(VIN), .Y(n37) );
  MX2X1 U18 ( .A(SR_to_MUL[29]), .B(SR_to_MUL[37]), .S0(VIN), .Y(n23) );
  MX2X1 U15 ( .A(SR_to_MUL[5]), .B(SR_to_MUL[13]), .S0(VIN), .Y(n20) );
  MX2X1 U6 ( .A(SR_to_MUL[31]), .B(SR_to_MUL[39]), .S0(VIN), .Y(n11) );
  MX2X1 U44 ( .A(SR_to_MUL[41]), .B(SR_to_MUL[49]), .S0(VIN), .Y(n49) );
  MX2X1 U8 ( .A(SR_to_MUL[47]), .B(SR_to_MUL[55]), .S0(VIN), .Y(n13) );
  MX2X1 U7 ( .A(SR_to_MUL[39]), .B(SR_to_MUL[47]), .S0(VIN), .Y(n12) );
  MX2X1 U3 ( .A(SR_to_MUL[15]), .B(SR_to_MUL[23]), .S0(VIN), .Y(n9) );
  MX2X1 U55 ( .A(SR_SRI_bit_temp_out[2]), .B(SR_SRI_bit_temp_out[1]), .S0(VIN), 
        .Y(n60) );
  MX2X1 U54 ( .A(SR_SRI_bit_temp_out[3]), .B(SR_SRI_bit_temp_out[2]), .S0(VIN), 
        .Y(n59) );
  MX2X1 U52 ( .A(SR_SRI_bit_temp_out[5]), .B(SR_SRI_bit_temp_out[4]), .S0(VIN), 
        .Y(n57) );
  MX2X1 U56 ( .A(SR_SRI_bit_temp_out[1]), .B(SR_SRI_bit_temp_out[0]), .S0(VIN), 
        .Y(n61) );
  MX2X1 U51 ( .A(SR_to_MUX), .B(SR_SRI_bit_temp_out[5]), .S0(VIN), .Y(n56) );
  MX2X1 U53 ( .A(SR_SRI_bit_temp_out[4]), .B(SR_SRI_bit_temp_out[3]), .S0(VIN), 
        .Y(n58) );
  ADDFX1 ADD2_2_add_16_DP_OP_276_702_2_U2 ( .A(
        ADD2_2_add_16_DP_OP_276_702_2_n18), .B(
        ADD2_2_add_16_DP_OP_276_702_2_n50), .CI(
        ADD2_2_add_16_DP_OP_276_702_2_n2), .CO(
        ADD2_2_add_16_DP_OP_276_702_2_n1), .S(ADD_esteso_11__16_) );
  ADDFX1 ADD2_2_add_16_DP_OP_276_702_2_U3 ( .A(
        ADD2_2_add_16_DP_OP_276_702_2_n19), .B(
        ADD2_2_add_16_DP_OP_276_702_2_n20), .CI(
        ADD2_2_add_16_DP_OP_276_702_2_n3), .CO(
        ADD2_2_add_16_DP_OP_276_702_2_n2), .S(ADD_esteso_11__15_) );
  ADDFX1 ADD2_2_add_16_DP_OP_276_702_2_U4 ( .A(
        ADD2_2_add_16_DP_OP_276_702_2_n21), .B(
        ADD2_2_add_16_DP_OP_276_702_2_n22), .CI(
        ADD2_2_add_16_DP_OP_276_702_2_n4), .CO(
        ADD2_2_add_16_DP_OP_276_702_2_n3), .S(ADD_esteso_11__14_) );
  ADDFX1 ADD2_2_add_16_DP_OP_276_702_2_U5 ( .A(
        ADD2_2_add_16_DP_OP_276_702_2_n23), .B(
        ADD2_2_add_16_DP_OP_276_702_2_n24), .CI(
        ADD2_2_add_16_DP_OP_276_702_2_n5), .CO(
        ADD2_2_add_16_DP_OP_276_702_2_n4), .S(ADD_esteso_11__13_) );
  ADDFX1 ADD2_2_add_16_DP_OP_276_702_2_U6 ( .A(
        ADD2_2_add_16_DP_OP_276_702_2_n25), .B(
        ADD2_2_add_16_DP_OP_276_702_2_n26), .CI(
        ADD2_2_add_16_DP_OP_276_702_2_n6), .CO(
        ADD2_2_add_16_DP_OP_276_702_2_n5), .S(ADD_esteso_11__12_) );
  ADDFX1 ADD2_2_add_16_DP_OP_276_702_2_U7 ( .A(
        ADD2_2_add_16_DP_OP_276_702_2_n27), .B(
        ADD2_2_add_16_DP_OP_276_702_2_n28), .CI(
        ADD2_2_add_16_DP_OP_276_702_2_n7), .CO(
        ADD2_2_add_16_DP_OP_276_702_2_n6), .S(ADD_esteso_11__11_) );
  ADDFX1 ADD2_2_add_16_DP_OP_276_702_2_U8 ( .A(
        ADD2_2_add_16_DP_OP_276_702_2_n29), .B(
        ADD2_2_add_16_DP_OP_276_702_2_n30), .CI(
        ADD2_2_add_16_DP_OP_276_702_2_n8), .CO(
        ADD2_2_add_16_DP_OP_276_702_2_n7), .S(ADD_esteso_11__10_) );
  ADDFX1 ADD2_2_add_16_DP_OP_276_702_2_U9 ( .A(
        ADD2_2_add_16_DP_OP_276_702_2_n31), .B(
        ADD2_2_add_16_DP_OP_276_702_2_n32), .CI(
        ADD2_2_add_16_DP_OP_276_702_2_n9), .CO(
        ADD2_2_add_16_DP_OP_276_702_2_n8), .S(ADD_esteso_11__9_) );
  ADDFX1 ADD2_2_add_16_DP_OP_276_702_2_U10 ( .A(
        ADD2_2_add_16_DP_OP_276_702_2_n33), .B(
        ADD2_2_add_16_DP_OP_276_702_2_n34), .CI(
        ADD2_2_add_16_DP_OP_276_702_2_n10), .CO(
        ADD2_2_add_16_DP_OP_276_702_2_n9), .S(ADD_esteso_11__8_) );
  ADDFX1 ADD2_2_add_16_DP_OP_276_702_2_U11 ( .A(
        ADD2_2_add_16_DP_OP_276_702_2_n35), .B(
        ADD2_2_add_16_DP_OP_276_702_2_n36), .CI(
        ADD2_2_add_16_DP_OP_276_702_2_n11), .CO(
        ADD2_2_add_16_DP_OP_276_702_2_n10), .S(ADD_esteso_11__7_) );
  ADDFX1 ADD2_2_add_16_DP_OP_276_702_2_U12 ( .A(
        ADD2_2_add_16_DP_OP_276_702_2_n37), .B(
        ADD2_2_add_16_DP_OP_276_702_2_n38), .CI(
        ADD2_2_add_16_DP_OP_276_702_2_n12), .CO(
        ADD2_2_add_16_DP_OP_276_702_2_n11), .S(ADD_esteso_11__6_) );
  ADDFX1 ADD2_2_add_16_DP_OP_276_702_2_U13 ( .A(
        ADD2_2_add_16_DP_OP_276_702_2_n39), .B(
        ADD2_2_add_16_DP_OP_276_702_2_n40), .CI(
        ADD2_2_add_16_DP_OP_276_702_2_n13), .CO(
        ADD2_2_add_16_DP_OP_276_702_2_n12), .S(ADD_esteso_11__5_) );
  ADDFX1 ADD2_2_add_16_DP_OP_276_702_2_U14 ( .A(
        ADD2_2_add_16_DP_OP_276_702_2_n41), .B(
        ADD2_2_add_16_DP_OP_276_702_2_n42), .CI(
        ADD2_2_add_16_DP_OP_276_702_2_n14), .CO(
        ADD2_2_add_16_DP_OP_276_702_2_n13), .S(ADD_esteso_11__4_) );
  ADDFX1 ADD2_2_add_16_DP_OP_276_702_2_U15 ( .A(
        ADD2_2_add_16_DP_OP_276_702_2_n43), .B(
        ADD2_2_add_16_DP_OP_276_702_2_n44), .CI(
        ADD2_2_add_16_DP_OP_276_702_2_n15), .CO(
        ADD2_2_add_16_DP_OP_276_702_2_n14), .S(ADD_esteso_11__3_) );
  ADDFX1 ADD2_2_add_16_DP_OP_276_702_2_U16 ( .A(
        ADD2_2_add_16_DP_OP_276_702_2_n45), .B(
        ADD2_2_add_16_DP_OP_276_702_2_n46), .CI(
        ADD2_2_add_16_DP_OP_276_702_2_n16), .CO(
        ADD2_2_add_16_DP_OP_276_702_2_n15), .S(ADD_esteso_11__2_) );
  ADDFX1 ADD2_2_add_16_DP_OP_276_702_2_U17 ( .A(
        ADD2_2_add_16_DP_OP_276_702_2_n17), .B(ADD_esteso_6__1_), .CI(
        ADD2_2_add_16_DP_OP_276_702_2_n47), .CO(
        ADD2_2_add_16_DP_OP_276_702_2_n16), .S(ADD_esteso_11__1_) );
  ADDFX1 ADD2_2_add_16_DP_OP_276_702_2_U18 ( .A(ADD_esteso_5__0_), .B(
        ADD_esteso_4__0_), .CI(ADD_esteso_6__0_), .CO(
        ADD2_2_add_16_DP_OP_276_702_2_n17), .S(ADD_esteso_11__0_) );
  ADDHX1 ADD2_2_add_16_DP_OP_276_702_2_U33 ( .A(ADD_esteso_5__1_), .B(
        ADD_esteso_4__1_), .CO(ADD2_2_add_16_DP_OP_276_702_2_n46), .S(
        ADD2_2_add_16_DP_OP_276_702_2_n47) );
  ADDFX1 ADD2_2_add_16_DP_OP_276_702_2_U32 ( .A(ADD_esteso_6__2_), .B(
        ADD_esteso_5__2_), .CI(ADD_esteso_4__2_), .CO(
        ADD2_2_add_16_DP_OP_276_702_2_n44), .S(
        ADD2_2_add_16_DP_OP_276_702_2_n45) );
  ADDFX1 ADD2_2_add_16_DP_OP_276_702_2_U31 ( .A(ADD_esteso_6__3_), .B(
        ADD_esteso_5__3_), .CI(ADD_esteso_4__3_), .CO(
        ADD2_2_add_16_DP_OP_276_702_2_n42), .S(
        ADD2_2_add_16_DP_OP_276_702_2_n43) );
  ADDFX1 ADD2_2_add_16_DP_OP_276_702_2_U30 ( .A(ADD_esteso_6__4_), .B(
        ADD_esteso_5__4_), .CI(ADD_esteso_4__4_), .CO(
        ADD2_2_add_16_DP_OP_276_702_2_n40), .S(
        ADD2_2_add_16_DP_OP_276_702_2_n41) );
  ADDFX1 ADD2_2_add_16_DP_OP_276_702_2_U29 ( .A(ADD_esteso_6__5_), .B(
        ADD_esteso_5__5_), .CI(ADD_esteso_4__5_), .CO(
        ADD2_2_add_16_DP_OP_276_702_2_n38), .S(
        ADD2_2_add_16_DP_OP_276_702_2_n39) );
  ADDFX1 ADD2_2_add_16_DP_OP_276_702_2_U28 ( .A(ADD_esteso_6__6_), .B(
        ADD_esteso_5__6_), .CI(ADD_esteso_4__6_), .CO(
        ADD2_2_add_16_DP_OP_276_702_2_n36), .S(
        ADD2_2_add_16_DP_OP_276_702_2_n37) );
  ADDFX1 ADD2_2_add_16_DP_OP_276_702_2_U27 ( .A(ADD_esteso_6__7_), .B(
        ADD_esteso_5__7_), .CI(ADD_esteso_4__7_), .CO(
        ADD2_2_add_16_DP_OP_276_702_2_n34), .S(
        ADD2_2_add_16_DP_OP_276_702_2_n35) );
  ADDFX1 ADD2_2_add_16_DP_OP_276_702_2_U26 ( .A(ADD_esteso_6__8_), .B(
        ADD_esteso_5__8_), .CI(ADD_esteso_4__8_), .CO(
        ADD2_2_add_16_DP_OP_276_702_2_n32), .S(
        ADD2_2_add_16_DP_OP_276_702_2_n33) );
  ADDFX1 ADD2_2_add_16_DP_OP_276_702_2_U25 ( .A(ADD_esteso_6__9_), .B(
        ADD_esteso_5__9_), .CI(ADD_esteso_4__9_), .CO(
        ADD2_2_add_16_DP_OP_276_702_2_n30), .S(
        ADD2_2_add_16_DP_OP_276_702_2_n31) );
  ADDFX1 ADD2_2_add_16_DP_OP_276_702_2_U24 ( .A(ADD_esteso_6__10_), .B(
        ADD_esteso_5__10_), .CI(ADD_esteso_4__10_), .CO(
        ADD2_2_add_16_DP_OP_276_702_2_n28), .S(
        ADD2_2_add_16_DP_OP_276_702_2_n29) );
  ADDFX1 ADD2_2_add_16_DP_OP_276_702_2_U23 ( .A(ADD_esteso_6__11_), .B(
        ADD_esteso_5__11_), .CI(ADD_esteso_4__11_), .CO(
        ADD2_2_add_16_DP_OP_276_702_2_n26), .S(
        ADD2_2_add_16_DP_OP_276_702_2_n27) );
  ADDFX1 ADD2_2_add_16_DP_OP_276_702_2_U22 ( .A(ADD_esteso_6__12_), .B(
        ADD_esteso_5__12_), .CI(ADD_esteso_4__12_), .CO(
        ADD2_2_add_16_DP_OP_276_702_2_n24), .S(
        ADD2_2_add_16_DP_OP_276_702_2_n25) );
  ADDFX1 ADD2_2_add_16_DP_OP_276_702_2_U21 ( .A(ADD_esteso_6__13_), .B(
        ADD_esteso_5__13_), .CI(ADD_esteso_4__13_), .CO(
        ADD2_2_add_16_DP_OP_276_702_2_n22), .S(
        ADD2_2_add_16_DP_OP_276_702_2_n23) );
  ADDFX1 ADD2_2_add_16_DP_OP_276_702_2_U20 ( .A(ADD_esteso_6__14_), .B(
        ADD_esteso_5__14_), .CI(ADD_esteso_4__14_), .CO(
        ADD2_2_add_16_DP_OP_276_702_2_n20), .S(
        ADD2_2_add_16_DP_OP_276_702_2_n21) );
  ADDFX1 ADD2_2_add_16_DP_OP_276_702_2_U19 ( .A(
        ADD2_2_add_16_DP_OP_276_702_2_n49), .B(ADD_esteso_5__17_), .CI(
        ADD2_2_add_16_DP_OP_276_702_2_n48), .CO(
        ADD2_2_add_16_DP_OP_276_702_2_n18), .S(
        ADD2_2_add_16_DP_OP_276_702_2_n19) );
  ADDFX1 ADD2_1_add_16_DP_OP_277_5600_1_U2 ( .A(
        ADD2_1_add_16_DP_OP_277_5600_1_n19), .B(
        ADD2_1_add_16_DP_OP_277_5600_1_n18), .CI(
        ADD2_1_add_16_DP_OP_277_5600_1_n2), .CO(
        ADD2_1_add_16_DP_OP_277_5600_1_n1), .S(ADD_esteso_10__16_) );
  ADDFX1 ADD2_1_add_16_DP_OP_277_5600_1_U3 ( .A(
        ADD2_1_add_16_DP_OP_277_5600_1_n20), .B(
        ADD2_1_add_16_DP_OP_277_5600_1_n22), .CI(
        ADD2_1_add_16_DP_OP_277_5600_1_n3), .CO(
        ADD2_1_add_16_DP_OP_277_5600_1_n2), .S(ADD_esteso_10__15_) );
  ADDFX1 ADD2_1_add_16_DP_OP_277_5600_1_U4 ( .A(
        ADD2_1_add_16_DP_OP_277_5600_1_n23), .B(
        ADD2_1_add_16_DP_OP_277_5600_1_n25), .CI(
        ADD2_1_add_16_DP_OP_277_5600_1_n4), .CO(
        ADD2_1_add_16_DP_OP_277_5600_1_n3), .S(ADD_esteso_10__14_) );
  ADDFX1 ADD2_1_add_16_DP_OP_277_5600_1_U5 ( .A(
        ADD2_1_add_16_DP_OP_277_5600_1_n26), .B(
        ADD2_1_add_16_DP_OP_277_5600_1_n28), .CI(
        ADD2_1_add_16_DP_OP_277_5600_1_n5), .CO(
        ADD2_1_add_16_DP_OP_277_5600_1_n4), .S(ADD_esteso_10__13_) );
  ADDFX1 ADD2_1_add_16_DP_OP_277_5600_1_U6 ( .A(
        ADD2_1_add_16_DP_OP_277_5600_1_n29), .B(
        ADD2_1_add_16_DP_OP_277_5600_1_n31), .CI(
        ADD2_1_add_16_DP_OP_277_5600_1_n6), .CO(
        ADD2_1_add_16_DP_OP_277_5600_1_n5), .S(ADD_esteso_10__12_) );
  ADDFX1 ADD2_1_add_16_DP_OP_277_5600_1_U7 ( .A(
        ADD2_1_add_16_DP_OP_277_5600_1_n32), .B(
        ADD2_1_add_16_DP_OP_277_5600_1_n34), .CI(
        ADD2_1_add_16_DP_OP_277_5600_1_n7), .CO(
        ADD2_1_add_16_DP_OP_277_5600_1_n6), .S(ADD_esteso_10__11_) );
  ADDFX1 ADD2_1_add_16_DP_OP_277_5600_1_U8 ( .A(
        ADD2_1_add_16_DP_OP_277_5600_1_n35), .B(
        ADD2_1_add_16_DP_OP_277_5600_1_n37), .CI(
        ADD2_1_add_16_DP_OP_277_5600_1_n8), .CO(
        ADD2_1_add_16_DP_OP_277_5600_1_n7), .S(ADD_esteso_10__10_) );
  ADDFX1 ADD2_1_add_16_DP_OP_277_5600_1_U9 ( .A(
        ADD2_1_add_16_DP_OP_277_5600_1_n38), .B(
        ADD2_1_add_16_DP_OP_277_5600_1_n40), .CI(
        ADD2_1_add_16_DP_OP_277_5600_1_n9), .CO(
        ADD2_1_add_16_DP_OP_277_5600_1_n8), .S(ADD_esteso_10__9_) );
  ADDFX1 ADD2_1_add_16_DP_OP_277_5600_1_U10 ( .A(
        ADD2_1_add_16_DP_OP_277_5600_1_n41), .B(
        ADD2_1_add_16_DP_OP_277_5600_1_n43), .CI(
        ADD2_1_add_16_DP_OP_277_5600_1_n10), .CO(
        ADD2_1_add_16_DP_OP_277_5600_1_n9), .S(ADD_esteso_10__8_) );
  ADDFX1 ADD2_1_add_16_DP_OP_277_5600_1_U11 ( .A(
        ADD2_1_add_16_DP_OP_277_5600_1_n44), .B(
        ADD2_1_add_16_DP_OP_277_5600_1_n46), .CI(
        ADD2_1_add_16_DP_OP_277_5600_1_n11), .CO(
        ADD2_1_add_16_DP_OP_277_5600_1_n10), .S(ADD_esteso_10__7_) );
  ADDFX1 ADD2_1_add_16_DP_OP_277_5600_1_U12 ( .A(
        ADD2_1_add_16_DP_OP_277_5600_1_n47), .B(
        ADD2_1_add_16_DP_OP_277_5600_1_n49), .CI(
        ADD2_1_add_16_DP_OP_277_5600_1_n12), .CO(
        ADD2_1_add_16_DP_OP_277_5600_1_n11), .S(ADD_esteso_10__6_) );
  ADDFX1 ADD2_1_add_16_DP_OP_277_5600_1_U13 ( .A(
        ADD2_1_add_16_DP_OP_277_5600_1_n50), .B(
        ADD2_1_add_16_DP_OP_277_5600_1_n52), .CI(
        ADD2_1_add_16_DP_OP_277_5600_1_n13), .CO(
        ADD2_1_add_16_DP_OP_277_5600_1_n12), .S(ADD_esteso_10__5_) );
  ADDFX1 ADD2_1_add_16_DP_OP_277_5600_1_U14 ( .A(
        ADD2_1_add_16_DP_OP_277_5600_1_n53), .B(
        ADD2_1_add_16_DP_OP_277_5600_1_n55), .CI(
        ADD2_1_add_16_DP_OP_277_5600_1_n14), .CO(
        ADD2_1_add_16_DP_OP_277_5600_1_n13), .S(ADD_esteso_10__4_) );
  ADDFX1 ADD2_1_add_16_DP_OP_277_5600_1_U15 ( .A(
        ADD2_1_add_16_DP_OP_277_5600_1_n56), .B(
        ADD2_1_add_16_DP_OP_277_5600_1_n58), .CI(
        ADD2_1_add_16_DP_OP_277_5600_1_n15), .CO(
        ADD2_1_add_16_DP_OP_277_5600_1_n14), .S(ADD_esteso_10__3_) );
  ADDFX1 ADD2_1_add_16_DP_OP_277_5600_1_U16 ( .A(
        ADD2_1_add_16_DP_OP_277_5600_1_n59), .B(
        ADD2_1_add_16_DP_OP_277_5600_1_n60), .CI(
        ADD2_1_add_16_DP_OP_277_5600_1_n16), .CO(
        ADD2_1_add_16_DP_OP_277_5600_1_n15), .S(ADD_esteso_10__2_) );
  ADDFX1 ADD2_1_add_16_DP_OP_277_5600_1_U17 ( .A(
        ADD2_1_add_16_DP_OP_277_5600_1_n61), .B(
        ADD2_1_add_16_DP_OP_277_5600_1_n63), .CI(
        ADD2_1_add_16_DP_OP_277_5600_1_n17), .CO(
        ADD2_1_add_16_DP_OP_277_5600_1_n16), .S(ADD_esteso_10__1_) );
  ADDFX1 ADD2_1_add_16_DP_OP_277_5600_1_U18 ( .A(ADD_esteso_3__0_), .B(
        ADD_esteso_0__0_), .CI(ADD2_1_add_16_DP_OP_277_5600_1_n65), .CO(
        ADD2_1_add_16_DP_OP_277_5600_1_n17), .S(ADD_esteso_10__0_) );
  ADDHX1 ADD2_1_add_16_DP_OP_277_5600_1_U34 ( .A(ADD_esteso_1__1_), .B(
        ADD_esteso_3__1_), .CO(ADD2_1_add_16_DP_OP_277_5600_1_n62), .S(
        ADD2_1_add_16_DP_OP_277_5600_1_n63) );
  ADDFX1 ADD2_1_add_16_DP_OP_277_5600_1_U33 ( .A(ADD_esteso_0__1_), .B(
        ADD_esteso_2__1_), .CI(ADD2_1_add_16_DP_OP_277_5600_1_n64), .CO(
        ADD2_1_add_16_DP_OP_277_5600_1_n60), .S(
        ADD2_1_add_16_DP_OP_277_5600_1_n61) );
  ADDHX1 ADD2_1_add_16_DP_OP_277_5600_1_U35 ( .A(ADD_esteso_1__0_), .B(
        ADD_esteso_2__0_), .CO(ADD2_1_add_16_DP_OP_277_5600_1_n64), .S(
        ADD2_1_add_16_DP_OP_277_5600_1_n65) );
  CMPR42X1 ADD2_1_add_16_DP_OP_277_5600_1_U32 ( .A(ADD_esteso_1__2_), .B(
        ADD_esteso_3__2_), .C(ADD_esteso_0__2_), .D(ADD_esteso_2__2_), .ICI(
        ADD2_1_add_16_DP_OP_277_5600_1_n62), .S(
        ADD2_1_add_16_DP_OP_277_5600_1_n59), .ICO(
        ADD2_1_add_16_DP_OP_277_5600_1_n57), .CO(
        ADD2_1_add_16_DP_OP_277_5600_1_n58) );
  CMPR42X1 ADD2_1_add_16_DP_OP_277_5600_1_U31 ( .A(ADD_esteso_1__3_), .B(
        ADD_esteso_3__3_), .C(ADD_esteso_0__3_), .D(ADD_esteso_2__3_), .ICI(
        ADD2_1_add_16_DP_OP_277_5600_1_n57), .S(
        ADD2_1_add_16_DP_OP_277_5600_1_n56), .ICO(
        ADD2_1_add_16_DP_OP_277_5600_1_n54), .CO(
        ADD2_1_add_16_DP_OP_277_5600_1_n55) );
  CMPR42X1 ADD2_1_add_16_DP_OP_277_5600_1_U30 ( .A(ADD_esteso_1__4_), .B(
        ADD_esteso_3__4_), .C(ADD_esteso_0__4_), .D(ADD_esteso_2__4_), .ICI(
        ADD2_1_add_16_DP_OP_277_5600_1_n54), .S(
        ADD2_1_add_16_DP_OP_277_5600_1_n53), .ICO(
        ADD2_1_add_16_DP_OP_277_5600_1_n51), .CO(
        ADD2_1_add_16_DP_OP_277_5600_1_n52) );
  CMPR42X1 ADD2_1_add_16_DP_OP_277_5600_1_U29 ( .A(ADD_esteso_1__5_), .B(
        ADD_esteso_3__5_), .C(ADD_esteso_0__5_), .D(ADD_esteso_2__5_), .ICI(
        ADD2_1_add_16_DP_OP_277_5600_1_n51), .S(
        ADD2_1_add_16_DP_OP_277_5600_1_n50), .ICO(
        ADD2_1_add_16_DP_OP_277_5600_1_n48), .CO(
        ADD2_1_add_16_DP_OP_277_5600_1_n49) );
  CMPR42X1 ADD2_1_add_16_DP_OP_277_5600_1_U28 ( .A(ADD_esteso_1__6_), .B(
        ADD_esteso_3__6_), .C(ADD_esteso_0__6_), .D(ADD_esteso_2__6_), .ICI(
        ADD2_1_add_16_DP_OP_277_5600_1_n48), .S(
        ADD2_1_add_16_DP_OP_277_5600_1_n47), .ICO(
        ADD2_1_add_16_DP_OP_277_5600_1_n45), .CO(
        ADD2_1_add_16_DP_OP_277_5600_1_n46) );
  CMPR42X1 ADD2_1_add_16_DP_OP_277_5600_1_U27 ( .A(ADD_esteso_1__7_), .B(
        ADD_esteso_3__7_), .C(ADD_esteso_0__7_), .D(ADD_esteso_2__7_), .ICI(
        ADD2_1_add_16_DP_OP_277_5600_1_n45), .S(
        ADD2_1_add_16_DP_OP_277_5600_1_n44), .ICO(
        ADD2_1_add_16_DP_OP_277_5600_1_n42), .CO(
        ADD2_1_add_16_DP_OP_277_5600_1_n43) );
  CMPR42X1 ADD2_1_add_16_DP_OP_277_5600_1_U26 ( .A(ADD_esteso_1__8_), .B(
        ADD_esteso_3__8_), .C(ADD_esteso_0__8_), .D(ADD_esteso_2__8_), .ICI(
        ADD2_1_add_16_DP_OP_277_5600_1_n42), .S(
        ADD2_1_add_16_DP_OP_277_5600_1_n41), .ICO(
        ADD2_1_add_16_DP_OP_277_5600_1_n39), .CO(
        ADD2_1_add_16_DP_OP_277_5600_1_n40) );
  CMPR42X1 ADD2_1_add_16_DP_OP_277_5600_1_U25 ( .A(ADD_esteso_1__9_), .B(
        ADD_esteso_3__9_), .C(ADD_esteso_0__9_), .D(ADD_esteso_2__9_), .ICI(
        ADD2_1_add_16_DP_OP_277_5600_1_n39), .S(
        ADD2_1_add_16_DP_OP_277_5600_1_n38), .ICO(
        ADD2_1_add_16_DP_OP_277_5600_1_n36), .CO(
        ADD2_1_add_16_DP_OP_277_5600_1_n37) );
  CMPR42X1 ADD2_1_add_16_DP_OP_277_5600_1_U24 ( .A(ADD_esteso_1__10_), .B(
        ADD_esteso_3__10_), .C(ADD_esteso_0__10_), .D(ADD_esteso_2__10_), 
        .ICI(ADD2_1_add_16_DP_OP_277_5600_1_n36), .S(
        ADD2_1_add_16_DP_OP_277_5600_1_n35), .ICO(
        ADD2_1_add_16_DP_OP_277_5600_1_n33), .CO(
        ADD2_1_add_16_DP_OP_277_5600_1_n34) );
  CMPR42X1 ADD2_1_add_16_DP_OP_277_5600_1_U23 ( .A(ADD_esteso_1__11_), .B(
        ADD_esteso_3__11_), .C(ADD_esteso_0__11_), .D(ADD_esteso_2__11_), 
        .ICI(ADD2_1_add_16_DP_OP_277_5600_1_n33), .S(
        ADD2_1_add_16_DP_OP_277_5600_1_n32), .ICO(
        ADD2_1_add_16_DP_OP_277_5600_1_n30), .CO(
        ADD2_1_add_16_DP_OP_277_5600_1_n31) );
  CMPR42X1 ADD2_1_add_16_DP_OP_277_5600_1_U22 ( .A(ADD_esteso_1__12_), .B(
        ADD_esteso_3__12_), .C(ADD_esteso_0__12_), .D(ADD_esteso_2__12_), 
        .ICI(ADD2_1_add_16_DP_OP_277_5600_1_n30), .S(
        ADD2_1_add_16_DP_OP_277_5600_1_n29), .ICO(
        ADD2_1_add_16_DP_OP_277_5600_1_n27), .CO(
        ADD2_1_add_16_DP_OP_277_5600_1_n28) );
  CMPR42X1 ADD2_1_add_16_DP_OP_277_5600_1_U21 ( .A(ADD_esteso_1__13_), .B(
        ADD_esteso_3__13_), .C(ADD_esteso_0__13_), .D(ADD_esteso_2__13_), 
        .ICI(ADD2_1_add_16_DP_OP_277_5600_1_n27), .S(
        ADD2_1_add_16_DP_OP_277_5600_1_n26), .ICO(
        ADD2_1_add_16_DP_OP_277_5600_1_n24), .CO(
        ADD2_1_add_16_DP_OP_277_5600_1_n25) );
  CMPR42X1 ADD2_1_add_16_DP_OP_277_5600_1_U20 ( .A(ADD_esteso_1__14_), .B(
        ADD_esteso_3__14_), .C(ADD_esteso_0__14_), .D(ADD_esteso_2__14_), 
        .ICI(ADD2_1_add_16_DP_OP_277_5600_1_n24), .S(
        ADD2_1_add_16_DP_OP_277_5600_1_n23), .ICO(
        ADD2_1_add_16_DP_OP_277_5600_1_n21), .CO(
        ADD2_1_add_16_DP_OP_277_5600_1_n22) );
  CMPR42X1 ADD2_1_add_16_DP_OP_277_5600_1_U19 ( .A(
        ADD2_1_add_16_DP_OP_277_5600_1_n21), .B(
        ADD2_1_add_16_DP_OP_277_5600_1_n67), .C(
        ADD2_1_add_16_DP_OP_277_5600_1_n66), .D(
        ADD2_1_add_16_DP_OP_277_5600_1_n68), .ICI(
        ADD2_1_add_16_DP_OP_277_5600_1_n69), .S(
        ADD2_1_add_16_DP_OP_277_5600_1_n20), .ICO(
        ADD2_1_add_16_DP_OP_277_5600_1_n18), .CO(
        ADD2_1_add_16_DP_OP_277_5600_1_n19) );
  ADDFX1 ADD3_1_add_16_U1_10 ( .A(ADD_esteso_12__10_), .B(ADD_esteso_13__10_), 
        .CI(ADD3_1_add_16_carry_10_), .CO(ADD3_1_add_16_carry_11_), .S(
        ADD_esteso_14__10_) );
  ADDFX1 ADD3_1_add_16_U1_11 ( .A(ADD_esteso_12__11_), .B(ADD_esteso_13__11_), 
        .CI(ADD3_1_add_16_carry_11_), .CO(ADD3_1_add_16_carry_12_), .S(
        ADD_esteso_14__11_) );
  ADDFX1 ADD3_1_add_16_U1_12 ( .A(ADD_esteso_12__12_), .B(ADD_esteso_13__12_), 
        .CI(ADD3_1_add_16_carry_12_), .CO(ADD3_1_add_16_carry_13_), .S(
        ADD_esteso_14__12_) );
  ADDFX1 ADD3_1_add_16_U1_13 ( .A(ADD_esteso_12__13_), .B(ADD_esteso_13__13_), 
        .CI(ADD3_1_add_16_carry_13_), .CO(ADD3_1_add_16_carry_14_), .S(
        ADD_esteso_14__13_) );
  ADDFX1 ADD3_1_add_16_U1_17 ( .A(ADD_esteso_12__17_), .B(ADD_esteso_13__17_), 
        .CI(ADD3_1_add_16_carry_17_), .S(ADD_esteso_14__17_) );
  ADDFX1 ADD3_1_add_16_U1_14 ( .A(ADD_esteso_12__14_), .B(ADD_esteso_13__14_), 
        .CI(ADD3_1_add_16_carry_14_), .CO(ADD3_1_add_16_carry_15_), .S(
        ADD_esteso_14__14_) );
  ADDFX1 ADD3_1_add_16_U1_15 ( .A(ADD_esteso_12__15_), .B(ADD_esteso_13__15_), 
        .CI(ADD3_1_add_16_carry_15_), .CO(ADD3_1_add_16_carry_16_), .S(
        ADD_esteso_14__15_) );
  ADDFX1 ADD3_1_add_16_U1_16 ( .A(ADD_esteso_12__16_), .B(ADD_esteso_13__16_), 
        .CI(ADD3_1_add_16_carry_16_), .CO(ADD3_1_add_16_carry_17_), .S(
        ADD_esteso_14__16_) );
  ADDFX1 MULi_1_mult_15_U5 ( .A(MULi_1_mult_15_n24), .B(MULi_1_mult_15_n20), 
        .CI(MULi_1_mult_15_n5), .CO(MULi_1_mult_15_n4), .S(MUL_to_PIPE1[91])
         );
  ADDFX1 MULi_1_mult_15_U6 ( .A(MULi_1_mult_15_n27), .B(MULi_1_mult_15_n25), 
        .CI(MULi_1_mult_15_n6), .CO(MULi_1_mult_15_n5), .S(MUL_to_PIPE1[90])
         );
  ADDFX1 MULi_1_mult_15_U7 ( .A(MULi_1_mult_15_n28), .B(MULi_1_mult_15_n32), 
        .CI(MULi_1_mult_15_n7), .CO(MULi_1_mult_15_n6), .S(MUL_to_PIPE1[89])
         );
  ADDFX1 MULi_1_mult_15_U8 ( .A(MULi_1_mult_15_n33), .B(MULi_1_mult_15_n37), 
        .CI(MULi_1_mult_15_n8), .CO(MULi_1_mult_15_n7), .S(MUL_to_PIPE1[88])
         );
  ADDFX1 MULi_1_mult_15_U9 ( .A(MULi_1_mult_15_n38), .B(MULi_1_mult_15_n42), 
        .CI(MULi_1_mult_15_n9), .CO(MULi_1_mult_15_n8), .S(MUL_to_PIPE1[87])
         );
  ADDFX1 MULi_1_mult_15_U10 ( .A(MULi_1_mult_15_n44), .B(MULi_1_mult_15_n43), 
        .CI(MULi_1_mult_15_n10), .CO(MULi_1_mult_15_n9), .S(MUL_to_PIPE1[86])
         );
  ADDFX1 MULi_1_mult_15_U11 ( .A(MULi_1_mult_15_n45), .B(MULi_1_mult_15_n47), 
        .CI(MULi_1_mult_15_n11), .CO(MULi_1_mult_15_n10), .S(MUL_to_PIPE1[85])
         );
  ADDFX1 MULi_1_mult_15_U12 ( .A(MULi_1_mult_15_n49), .B(MULi_1_mult_15_n50), 
        .CI(MULi_1_mult_15_n12), .CO(MULi_1_mult_15_n11), .S(MUL_to_PIPE1[84])
         );
  ADDFX1 MULi_1_mult_15_U13 ( .A(MULi_1_mult_15_n51), .B(MULi_1_mult_15_n54), 
        .CI(MULi_1_mult_15_n13), .CO(MULi_1_mult_15_n12), .S(MUL_to_PIPE1[83])
         );
  ADDFX1 MULi_1_mult_15_U14 ( .A(MULi_1_mult_15_n86), .B(MULi_1_mult_15_n79), 
        .CI(MULi_1_mult_15_n14), .CO(MULi_1_mult_15_n13), .S(MUL_to_PIPE1[82])
         );
  ADDHX1 MULi_1_mult_15_U15 ( .A(MULi_1_mult_15_n55), .B(MULi_1_mult_15_n87), 
        .CO(MULi_1_mult_15_n14), .S(MUL_to_PIPE1[81]) );
  ADDFX1 MULi_1_mult_15_U29 ( .A(MULi_1_mult_15_n70), .B(MULi_1_mult_15_n76), 
        .CI(MULi_1_mult_15_n48), .CO(MULi_1_mult_15_n44), .S(
        MULi_1_mult_15_n45) );
  ADDFX1 MULi_1_mult_15_U31 ( .A(MULi_1_mult_15_n84), .B(MULi_1_mult_15_n71), 
        .CI(MULi_1_mult_15_n77), .CO(MULi_1_mult_15_n48), .S(
        MULi_1_mult_15_n49) );
  ADDFX1 MULi_1_mult_15_U18 ( .A(MULi_1_mult_15_n22), .B(MULi_1_mult_15_n58), 
        .CI(MULi_1_mult_15_n23), .CO(MULi_1_mult_15_n19), .S(
        MULi_1_mult_15_n20) );
  ADDFX1 MULi_1_mult_15_U17 ( .A(MULi_1_mult_15_n57), .B(MULi_1_mult_15_n64), 
        .CI(MULi_1_mult_15_n21), .CO(MULi_1_mult_15_n17), .S(
        MULi_1_mult_15_n18) );
  CMPR42X1 MULi_1_mult_15_U28 ( .A(MULi_1_mult_15_n63), .B(MULi_1_mult_15_n82), 
        .C(MULi_1_mult_15_n75), .D(MULi_1_mult_15_n69), .ICI(
        MULi_1_mult_15_n46), .S(MULi_1_mult_15_n43), .ICO(MULi_1_mult_15_n41), 
        .CO(MULi_1_mult_15_n42) );
  CMPR42X1 MULi_1_mult_15_U26 ( .A(MULi_1_mult_15_n74), .B(MULi_1_mult_15_n62), 
        .C(MULi_1_mult_15_n68), .D(MULi_1_mult_15_n41), .ICI(
        MULi_1_mult_15_n40), .S(MULi_1_mult_15_n38), .ICO(MULi_1_mult_15_n36), 
        .CO(MULi_1_mult_15_n37) );
  CMPR42X1 MULi_1_mult_15_U23 ( .A(MULi_1_mult_15_n67), .B(MULi_1_mult_15_n61), 
        .C(MULi_1_mult_15_n39), .D(MULi_1_mult_15_n36), .ICI(
        MULi_1_mult_15_n35), .S(MULi_1_mult_15_n33), .ICO(MULi_1_mult_15_n31), 
        .CO(MULi_1_mult_15_n32) );
  CMPR42X1 MULi_1_mult_15_U21 ( .A(MULi_1_mult_15_n66), .B(MULi_1_mult_15_n60), 
        .C(n169), .D(MULi_1_mult_15_n34), .ICI(MULi_1_mult_15_n31), .S(
        MULi_1_mult_15_n28), .ICO(MULi_1_mult_15_n26), .CO(MULi_1_mult_15_n27)
         );
  CMPR42X1 MULi_1_mult_15_U20 ( .A(MULi_1_mult_15_n72), .B(MULi_1_mult_15_n65), 
        .C(MULi_1_mult_15_n59), .D(n168), .ICI(MULi_1_mult_15_n26), .S(
        MULi_1_mult_15_n25), .ICO(MULi_1_mult_15_n23), .CO(MULi_1_mult_15_n24)
         );
  ADDFX1 MULi_2_mult_15_U2 ( .A(MULi_2_mult_15_n15), .B(MULi_2_mult_15_n56), 
        .CI(MULi_2_mult_15_n2), .CO(MULi_2_mult_15_n1), .S(MUL_to_PIPE1[78])
         );
  ADDFX1 MULi_2_mult_15_U3 ( .A(MULi_2_mult_15_n17), .B(MULi_2_mult_15_n16), 
        .CI(MULi_2_mult_15_n3), .CO(MULi_2_mult_15_n2), .S(MUL_to_PIPE1[77])
         );
  ADDFX1 MULi_2_mult_15_U4 ( .A(MULi_2_mult_15_n19), .B(MULi_2_mult_15_n18), 
        .CI(MULi_2_mult_15_n4), .CO(MULi_2_mult_15_n3), .S(MUL_to_PIPE1[76])
         );
  ADDFX1 MULi_2_mult_15_U5 ( .A(MULi_2_mult_15_n24), .B(MULi_2_mult_15_n20), 
        .CI(MULi_2_mult_15_n5), .CO(MULi_2_mult_15_n4), .S(MUL_to_PIPE1[75])
         );
  ADDFX1 MULi_2_mult_15_U6 ( .A(MULi_2_mult_15_n27), .B(MULi_2_mult_15_n25), 
        .CI(MULi_2_mult_15_n6), .CO(MULi_2_mult_15_n5), .S(MUL_to_PIPE1[74])
         );
  ADDFX1 MULi_2_mult_15_U7 ( .A(MULi_2_mult_15_n28), .B(MULi_2_mult_15_n32), 
        .CI(MULi_2_mult_15_n7), .CO(MULi_2_mult_15_n6), .S(MUL_to_PIPE1[73])
         );
  ADDFX1 MULi_2_mult_15_U8 ( .A(MULi_2_mult_15_n33), .B(MULi_2_mult_15_n37), 
        .CI(MULi_2_mult_15_n8), .CO(MULi_2_mult_15_n7), .S(MUL_to_PIPE1[72])
         );
  ADDFX1 MULi_2_mult_15_U9 ( .A(MULi_2_mult_15_n38), .B(MULi_2_mult_15_n42), 
        .CI(MULi_2_mult_15_n9), .CO(MULi_2_mult_15_n8), .S(MUL_to_PIPE1[71])
         );
  ADDFX1 MULi_2_mult_15_U10 ( .A(MULi_2_mult_15_n44), .B(MULi_2_mult_15_n43), 
        .CI(MULi_2_mult_15_n10), .CO(MULi_2_mult_15_n9), .S(MUL_to_PIPE1[70])
         );
  ADDFX1 MULi_2_mult_15_U11 ( .A(MULi_2_mult_15_n45), .B(MULi_2_mult_15_n47), 
        .CI(MULi_2_mult_15_n11), .CO(MULi_2_mult_15_n10), .S(MUL_to_PIPE1[69])
         );
  ADDFX1 MULi_2_mult_15_U12 ( .A(MULi_2_mult_15_n49), .B(MULi_2_mult_15_n50), 
        .CI(MULi_2_mult_15_n12), .CO(MULi_2_mult_15_n11), .S(MUL_to_PIPE1[68])
         );
  ADDFX1 MULi_2_mult_15_U13 ( .A(MULi_2_mult_15_n51), .B(MULi_2_mult_15_n54), 
        .CI(MULi_2_mult_15_n13), .CO(MULi_2_mult_15_n12), .S(MUL_to_PIPE1[67])
         );
  ADDFX1 MULi_2_mult_15_U14 ( .A(MULi_2_mult_15_n86), .B(MULi_2_mult_15_n79), 
        .CI(MULi_2_mult_15_n14), .CO(MULi_2_mult_15_n13), .S(MUL_to_PIPE1[66])
         );
  ADDHX1 MULi_2_mult_15_U15 ( .A(MULi_2_mult_15_n55), .B(MULi_2_mult_15_n87), 
        .CO(MULi_2_mult_15_n14), .S(MUL_to_PIPE1[65]) );
  ADDFX1 MULi_2_mult_15_U29 ( .A(MULi_2_mult_15_n70), .B(MULi_2_mult_15_n76), 
        .CI(MULi_2_mult_15_n48), .CO(MULi_2_mult_15_n44), .S(
        MULi_2_mult_15_n45) );
  ADDFX1 MULi_2_mult_15_U31 ( .A(MULi_2_mult_15_n84), .B(MULi_2_mult_15_n71), 
        .CI(MULi_2_mult_15_n77), .CO(MULi_2_mult_15_n48), .S(
        MULi_2_mult_15_n49) );
  ADDFX1 MULi_2_mult_15_U18 ( .A(MULi_2_mult_15_n22), .B(MULi_2_mult_15_n58), 
        .CI(MULi_2_mult_15_n23), .CO(MULi_2_mult_15_n19), .S(
        MULi_2_mult_15_n20) );
  ADDFX1 MULi_2_mult_15_U17 ( .A(MULi_2_mult_15_n57), .B(MULi_2_mult_15_n64), 
        .CI(MULi_2_mult_15_n21), .CO(MULi_2_mult_15_n17), .S(
        MULi_2_mult_15_n18) );
  CMPR42X1 MULi_2_mult_15_U28 ( .A(MULi_2_mult_15_n63), .B(MULi_2_mult_15_n82), 
        .C(MULi_2_mult_15_n75), .D(MULi_2_mult_15_n69), .ICI(
        MULi_2_mult_15_n46), .S(MULi_2_mult_15_n43), .ICO(MULi_2_mult_15_n41), 
        .CO(MULi_2_mult_15_n42) );
  CMPR42X1 MULi_2_mult_15_U26 ( .A(MULi_2_mult_15_n74), .B(MULi_2_mult_15_n62), 
        .C(MULi_2_mult_15_n68), .D(MULi_2_mult_15_n41), .ICI(
        MULi_2_mult_15_n40), .S(MULi_2_mult_15_n38), .ICO(MULi_2_mult_15_n36), 
        .CO(MULi_2_mult_15_n37) );
  CMPR42X1 MULi_2_mult_15_U23 ( .A(MULi_2_mult_15_n67), .B(MULi_2_mult_15_n61), 
        .C(MULi_2_mult_15_n39), .D(MULi_2_mult_15_n36), .ICI(
        MULi_2_mult_15_n35), .S(MULi_2_mult_15_n33), .ICO(MULi_2_mult_15_n31), 
        .CO(MULi_2_mult_15_n32) );
  CMPR42X1 MULi_2_mult_15_U21 ( .A(MULi_2_mult_15_n66), .B(MULi_2_mult_15_n60), 
        .C(n165), .D(MULi_2_mult_15_n34), .ICI(MULi_2_mult_15_n31), .S(
        MULi_2_mult_15_n28), .ICO(MULi_2_mult_15_n26), .CO(MULi_2_mult_15_n27)
         );
  CMPR42X1 MULi_2_mult_15_U20 ( .A(MULi_2_mult_15_n72), .B(MULi_2_mult_15_n65), 
        .C(MULi_2_mult_15_n59), .D(n164), .ICI(MULi_2_mult_15_n26), .S(
        MULi_2_mult_15_n25), .ICO(MULi_2_mult_15_n23), .CO(MULi_2_mult_15_n24)
         );
  ADDFX1 MULi_3_mult_15_U5 ( .A(MULi_3_mult_15_n24), .B(MULi_3_mult_15_n20), 
        .CI(MULi_3_mult_15_n5), .CO(MULi_3_mult_15_n4), .S(MUL_to_PIPE1[59])
         );
  ADDFX1 MULi_3_mult_15_U6 ( .A(MULi_3_mult_15_n27), .B(MULi_3_mult_15_n25), 
        .CI(MULi_3_mult_15_n6), .CO(MULi_3_mult_15_n5), .S(MUL_to_PIPE1[58])
         );
  ADDFX1 MULi_3_mult_15_U7 ( .A(MULi_3_mult_15_n28), .B(MULi_3_mult_15_n32), 
        .CI(MULi_3_mult_15_n7), .CO(MULi_3_mult_15_n6), .S(MUL_to_PIPE1[57])
         );
  ADDFX1 MULi_3_mult_15_U8 ( .A(MULi_3_mult_15_n33), .B(MULi_3_mult_15_n37), 
        .CI(MULi_3_mult_15_n8), .CO(MULi_3_mult_15_n7), .S(MUL_to_PIPE1[56])
         );
  ADDFX1 MULi_3_mult_15_U9 ( .A(MULi_3_mult_15_n38), .B(MULi_3_mult_15_n42), 
        .CI(MULi_3_mult_15_n9), .CO(MULi_3_mult_15_n8), .S(MUL_to_PIPE1[55])
         );
  ADDFX1 MULi_3_mult_15_U10 ( .A(MULi_3_mult_15_n44), .B(MULi_3_mult_15_n43), 
        .CI(MULi_3_mult_15_n10), .CO(MULi_3_mult_15_n9), .S(MUL_to_PIPE1[54])
         );
  ADDFX1 MULi_3_mult_15_U11 ( .A(MULi_3_mult_15_n45), .B(MULi_3_mult_15_n47), 
        .CI(MULi_3_mult_15_n11), .CO(MULi_3_mult_15_n10), .S(MUL_to_PIPE1[53])
         );
  ADDFX1 MULi_3_mult_15_U12 ( .A(MULi_3_mult_15_n49), .B(MULi_3_mult_15_n50), 
        .CI(MULi_3_mult_15_n12), .CO(MULi_3_mult_15_n11), .S(MUL_to_PIPE1[52])
         );
  ADDFX1 MULi_3_mult_15_U13 ( .A(MULi_3_mult_15_n51), .B(MULi_3_mult_15_n54), 
        .CI(MULi_3_mult_15_n13), .CO(MULi_3_mult_15_n12), .S(MUL_to_PIPE1[51])
         );
  ADDFX1 MULi_3_mult_15_U14 ( .A(MULi_3_mult_15_n86), .B(MULi_3_mult_15_n79), 
        .CI(MULi_3_mult_15_n14), .CO(MULi_3_mult_15_n13), .S(MUL_to_PIPE1[50])
         );
  ADDHX1 MULi_3_mult_15_U15 ( .A(MULi_3_mult_15_n55), .B(MULi_3_mult_15_n87), 
        .CO(MULi_3_mult_15_n14), .S(MUL_to_PIPE1[49]) );
  ADDFX1 MULi_3_mult_15_U29 ( .A(MULi_3_mult_15_n70), .B(MULi_3_mult_15_n76), 
        .CI(MULi_3_mult_15_n48), .CO(MULi_3_mult_15_n44), .S(
        MULi_3_mult_15_n45) );
  ADDFX1 MULi_3_mult_15_U31 ( .A(MULi_3_mult_15_n84), .B(MULi_3_mult_15_n71), 
        .CI(MULi_3_mult_15_n77), .CO(MULi_3_mult_15_n48), .S(
        MULi_3_mult_15_n49) );
  ADDFX1 MULi_3_mult_15_U18 ( .A(MULi_3_mult_15_n22), .B(MULi_3_mult_15_n58), 
        .CI(MULi_3_mult_15_n23), .CO(MULi_3_mult_15_n19), .S(
        MULi_3_mult_15_n20) );
  ADDFX1 MULi_3_mult_15_U17 ( .A(MULi_3_mult_15_n57), .B(MULi_3_mult_15_n64), 
        .CI(MULi_3_mult_15_n21), .CO(MULi_3_mult_15_n17), .S(
        MULi_3_mult_15_n18) );
  CMPR42X1 MULi_3_mult_15_U28 ( .A(MULi_3_mult_15_n63), .B(MULi_3_mult_15_n82), 
        .C(MULi_3_mult_15_n75), .D(MULi_3_mult_15_n69), .ICI(
        MULi_3_mult_15_n46), .S(MULi_3_mult_15_n43), .ICO(MULi_3_mult_15_n41), 
        .CO(MULi_3_mult_15_n42) );
  CMPR42X1 MULi_3_mult_15_U26 ( .A(MULi_3_mult_15_n74), .B(MULi_3_mult_15_n62), 
        .C(MULi_3_mult_15_n68), .D(MULi_3_mult_15_n41), .ICI(
        MULi_3_mult_15_n40), .S(MULi_3_mult_15_n38), .ICO(MULi_3_mult_15_n36), 
        .CO(MULi_3_mult_15_n37) );
  CMPR42X1 MULi_3_mult_15_U23 ( .A(MULi_3_mult_15_n67), .B(MULi_3_mult_15_n61), 
        .C(MULi_3_mult_15_n39), .D(MULi_3_mult_15_n36), .ICI(
        MULi_3_mult_15_n35), .S(MULi_3_mult_15_n33), .ICO(MULi_3_mult_15_n31), 
        .CO(MULi_3_mult_15_n32) );
  CMPR42X1 MULi_3_mult_15_U21 ( .A(MULi_3_mult_15_n66), .B(MULi_3_mult_15_n60), 
        .C(n161), .D(MULi_3_mult_15_n34), .ICI(MULi_3_mult_15_n31), .S(
        MULi_3_mult_15_n28), .ICO(MULi_3_mult_15_n26), .CO(MULi_3_mult_15_n27)
         );
  CMPR42X1 MULi_3_mult_15_U20 ( .A(MULi_3_mult_15_n72), .B(MULi_3_mult_15_n65), 
        .C(MULi_3_mult_15_n59), .D(n160), .ICI(MULi_3_mult_15_n26), .S(
        MULi_3_mult_15_n25), .ICO(MULi_3_mult_15_n23), .CO(MULi_3_mult_15_n24)
         );
  ADDFX1 MULi_4_mult_15_U2 ( .A(MULi_4_mult_15_n15), .B(MULi_4_mult_15_n56), 
        .CI(MULi_4_mult_15_n2), .CO(MULi_4_mult_15_n1), .S(MUL_to_PIPE1[46])
         );
  ADDFX1 MULi_4_mult_15_U3 ( .A(MULi_4_mult_15_n17), .B(MULi_4_mult_15_n16), 
        .CI(MULi_4_mult_15_n3), .CO(MULi_4_mult_15_n2), .S(MUL_to_PIPE1[45])
         );
  ADDFX1 MULi_4_mult_15_U4 ( .A(MULi_4_mult_15_n19), .B(MULi_4_mult_15_n18), 
        .CI(MULi_4_mult_15_n4), .CO(MULi_4_mult_15_n3), .S(MUL_to_PIPE1[44])
         );
  ADDFX1 MULi_4_mult_15_U5 ( .A(MULi_4_mult_15_n24), .B(MULi_4_mult_15_n20), 
        .CI(MULi_4_mult_15_n5), .CO(MULi_4_mult_15_n4), .S(MUL_to_PIPE1[43])
         );
  ADDFX1 MULi_4_mult_15_U6 ( .A(MULi_4_mult_15_n27), .B(MULi_4_mult_15_n25), 
        .CI(MULi_4_mult_15_n6), .CO(MULi_4_mult_15_n5), .S(MUL_to_PIPE1[42])
         );
  ADDFX1 MULi_4_mult_15_U7 ( .A(MULi_4_mult_15_n28), .B(MULi_4_mult_15_n32), 
        .CI(MULi_4_mult_15_n7), .CO(MULi_4_mult_15_n6), .S(MUL_to_PIPE1[41])
         );
  ADDFX1 MULi_4_mult_15_U8 ( .A(MULi_4_mult_15_n33), .B(MULi_4_mult_15_n37), 
        .CI(MULi_4_mult_15_n8), .CO(MULi_4_mult_15_n7), .S(MUL_to_PIPE1[40])
         );
  ADDFX1 MULi_4_mult_15_U9 ( .A(MULi_4_mult_15_n38), .B(MULi_4_mult_15_n42), 
        .CI(MULi_4_mult_15_n9), .CO(MULi_4_mult_15_n8), .S(MUL_to_PIPE1[39])
         );
  ADDFX1 MULi_4_mult_15_U10 ( .A(MULi_4_mult_15_n44), .B(MULi_4_mult_15_n43), 
        .CI(MULi_4_mult_15_n10), .CO(MULi_4_mult_15_n9), .S(MUL_to_PIPE1[38])
         );
  ADDFX1 MULi_4_mult_15_U11 ( .A(MULi_4_mult_15_n45), .B(MULi_4_mult_15_n47), 
        .CI(MULi_4_mult_15_n11), .CO(MULi_4_mult_15_n10), .S(MUL_to_PIPE1[37])
         );
  ADDFX1 MULi_4_mult_15_U12 ( .A(MULi_4_mult_15_n49), .B(MULi_4_mult_15_n50), 
        .CI(MULi_4_mult_15_n12), .CO(MULi_4_mult_15_n11), .S(MUL_to_PIPE1[36])
         );
  ADDFX1 MULi_4_mult_15_U13 ( .A(MULi_4_mult_15_n51), .B(MULi_4_mult_15_n54), 
        .CI(MULi_4_mult_15_n13), .CO(MULi_4_mult_15_n12), .S(MUL_to_PIPE1[35])
         );
  ADDFX1 MULi_4_mult_15_U14 ( .A(MULi_4_mult_15_n86), .B(MULi_4_mult_15_n79), 
        .CI(MULi_4_mult_15_n14), .CO(MULi_4_mult_15_n13), .S(MUL_to_PIPE1[34])
         );
  ADDHX1 MULi_4_mult_15_U15 ( .A(MULi_4_mult_15_n55), .B(MULi_4_mult_15_n87), 
        .CO(MULi_4_mult_15_n14), .S(MUL_to_PIPE1[33]) );
  ADDFX1 MULi_4_mult_15_U29 ( .A(MULi_4_mult_15_n70), .B(MULi_4_mult_15_n76), 
        .CI(MULi_4_mult_15_n48), .CO(MULi_4_mult_15_n44), .S(
        MULi_4_mult_15_n45) );
  ADDFX1 MULi_4_mult_15_U31 ( .A(MULi_4_mult_15_n84), .B(MULi_4_mult_15_n71), 
        .CI(MULi_4_mult_15_n77), .CO(MULi_4_mult_15_n48), .S(
        MULi_4_mult_15_n49) );
  ADDFX1 MULi_4_mult_15_U18 ( .A(MULi_4_mult_15_n22), .B(MULi_4_mult_15_n58), 
        .CI(MULi_4_mult_15_n23), .CO(MULi_4_mult_15_n19), .S(
        MULi_4_mult_15_n20) );
  ADDFX1 MULi_4_mult_15_U17 ( .A(MULi_4_mult_15_n57), .B(MULi_4_mult_15_n64), 
        .CI(MULi_4_mult_15_n21), .CO(MULi_4_mult_15_n17), .S(
        MULi_4_mult_15_n18) );
  CMPR42X1 MULi_4_mult_15_U28 ( .A(MULi_4_mult_15_n63), .B(MULi_4_mult_15_n82), 
        .C(MULi_4_mult_15_n75), .D(MULi_4_mult_15_n69), .ICI(
        MULi_4_mult_15_n46), .S(MULi_4_mult_15_n43), .ICO(MULi_4_mult_15_n41), 
        .CO(MULi_4_mult_15_n42) );
  CMPR42X1 MULi_4_mult_15_U26 ( .A(MULi_4_mult_15_n74), .B(MULi_4_mult_15_n62), 
        .C(MULi_4_mult_15_n68), .D(MULi_4_mult_15_n41), .ICI(
        MULi_4_mult_15_n40), .S(MULi_4_mult_15_n38), .ICO(MULi_4_mult_15_n36), 
        .CO(MULi_4_mult_15_n37) );
  CMPR42X1 MULi_4_mult_15_U23 ( .A(MULi_4_mult_15_n67), .B(MULi_4_mult_15_n61), 
        .C(MULi_4_mult_15_n39), .D(MULi_4_mult_15_n36), .ICI(
        MULi_4_mult_15_n35), .S(MULi_4_mult_15_n33), .ICO(MULi_4_mult_15_n31), 
        .CO(MULi_4_mult_15_n32) );
  CMPR42X1 MULi_4_mult_15_U21 ( .A(MULi_4_mult_15_n66), .B(MULi_4_mult_15_n60), 
        .C(n159), .D(MULi_4_mult_15_n34), .ICI(MULi_4_mult_15_n31), .S(
        MULi_4_mult_15_n28), .ICO(MULi_4_mult_15_n26), .CO(MULi_4_mult_15_n27)
         );
  CMPR42X1 MULi_4_mult_15_U20 ( .A(MULi_4_mult_15_n72), .B(MULi_4_mult_15_n65), 
        .C(MULi_4_mult_15_n59), .D(n158), .ICI(MULi_4_mult_15_n26), .S(
        MULi_4_mult_15_n25), .ICO(MULi_4_mult_15_n23), .CO(MULi_4_mult_15_n24)
         );
  ADDFX1 MULi_5_mult_15_U5 ( .A(MULi_5_mult_15_n24), .B(MULi_5_mult_15_n20), 
        .CI(MULi_5_mult_15_n5), .CO(MULi_5_mult_15_n4), .S(MUL_to_PIPE1[27])
         );
  ADDFX1 MULi_5_mult_15_U6 ( .A(MULi_5_mult_15_n27), .B(MULi_5_mult_15_n25), 
        .CI(MULi_5_mult_15_n6), .CO(MULi_5_mult_15_n5), .S(MUL_to_PIPE1[26])
         );
  ADDFX1 MULi_5_mult_15_U7 ( .A(MULi_5_mult_15_n28), .B(MULi_5_mult_15_n32), 
        .CI(MULi_5_mult_15_n7), .CO(MULi_5_mult_15_n6), .S(MUL_to_PIPE1[25])
         );
  ADDFX1 MULi_5_mult_15_U8 ( .A(MULi_5_mult_15_n33), .B(MULi_5_mult_15_n37), 
        .CI(MULi_5_mult_15_n8), .CO(MULi_5_mult_15_n7), .S(MUL_to_PIPE1[24])
         );
  ADDFX1 MULi_5_mult_15_U9 ( .A(MULi_5_mult_15_n38), .B(MULi_5_mult_15_n42), 
        .CI(MULi_5_mult_15_n9), .CO(MULi_5_mult_15_n8), .S(MUL_to_PIPE1[23])
         );
  ADDFX1 MULi_5_mult_15_U10 ( .A(MULi_5_mult_15_n44), .B(MULi_5_mult_15_n43), 
        .CI(MULi_5_mult_15_n10), .CO(MULi_5_mult_15_n9), .S(MUL_to_PIPE1[22])
         );
  ADDFX1 MULi_5_mult_15_U11 ( .A(MULi_5_mult_15_n45), .B(MULi_5_mult_15_n47), 
        .CI(MULi_5_mult_15_n11), .CO(MULi_5_mult_15_n10), .S(MUL_to_PIPE1[21])
         );
  ADDFX1 MULi_5_mult_15_U12 ( .A(MULi_5_mult_15_n49), .B(MULi_5_mult_15_n50), 
        .CI(MULi_5_mult_15_n12), .CO(MULi_5_mult_15_n11), .S(MUL_to_PIPE1[20])
         );
  ADDFX1 MULi_5_mult_15_U13 ( .A(MULi_5_mult_15_n51), .B(MULi_5_mult_15_n54), 
        .CI(MULi_5_mult_15_n13), .CO(MULi_5_mult_15_n12), .S(MUL_to_PIPE1[19])
         );
  ADDFX1 MULi_5_mult_15_U14 ( .A(MULi_5_mult_15_n86), .B(MULi_5_mult_15_n79), 
        .CI(MULi_5_mult_15_n14), .CO(MULi_5_mult_15_n13), .S(MUL_to_PIPE1[18])
         );
  ADDHX1 MULi_5_mult_15_U15 ( .A(MULi_5_mult_15_n55), .B(MULi_5_mult_15_n87), 
        .CO(MULi_5_mult_15_n14), .S(MUL_to_PIPE1[17]) );
  ADDFX1 MULi_5_mult_15_U29 ( .A(MULi_5_mult_15_n70), .B(MULi_5_mult_15_n76), 
        .CI(MULi_5_mult_15_n48), .CO(MULi_5_mult_15_n44), .S(
        MULi_5_mult_15_n45) );
  ADDFX1 MULi_5_mult_15_U31 ( .A(MULi_5_mult_15_n84), .B(MULi_5_mult_15_n71), 
        .CI(MULi_5_mult_15_n77), .CO(MULi_5_mult_15_n48), .S(
        MULi_5_mult_15_n49) );
  ADDFX1 MULi_5_mult_15_U18 ( .A(MULi_5_mult_15_n22), .B(MULi_5_mult_15_n58), 
        .CI(MULi_5_mult_15_n23), .CO(MULi_5_mult_15_n19), .S(
        MULi_5_mult_15_n20) );
  ADDFX1 MULi_5_mult_15_U17 ( .A(MULi_5_mult_15_n57), .B(MULi_5_mult_15_n64), 
        .CI(MULi_5_mult_15_n21), .CO(MULi_5_mult_15_n17), .S(
        MULi_5_mult_15_n18) );
  CMPR42X1 MULi_5_mult_15_U28 ( .A(MULi_5_mult_15_n63), .B(MULi_5_mult_15_n82), 
        .C(MULi_5_mult_15_n75), .D(MULi_5_mult_15_n69), .ICI(
        MULi_5_mult_15_n46), .S(MULi_5_mult_15_n43), .ICO(MULi_5_mult_15_n41), 
        .CO(MULi_5_mult_15_n42) );
  CMPR42X1 MULi_5_mult_15_U26 ( .A(MULi_5_mult_15_n74), .B(MULi_5_mult_15_n62), 
        .C(MULi_5_mult_15_n68), .D(MULi_5_mult_15_n41), .ICI(
        MULi_5_mult_15_n40), .S(MULi_5_mult_15_n38), .ICO(MULi_5_mult_15_n36), 
        .CO(MULi_5_mult_15_n37) );
  CMPR42X1 MULi_5_mult_15_U23 ( .A(MULi_5_mult_15_n67), .B(MULi_5_mult_15_n61), 
        .C(MULi_5_mult_15_n39), .D(MULi_5_mult_15_n36), .ICI(
        MULi_5_mult_15_n35), .S(MULi_5_mult_15_n33), .ICO(MULi_5_mult_15_n31), 
        .CO(MULi_5_mult_15_n32) );
  CMPR42X1 MULi_5_mult_15_U21 ( .A(MULi_5_mult_15_n66), .B(MULi_5_mult_15_n60), 
        .C(n163), .D(MULi_5_mult_15_n34), .ICI(MULi_5_mult_15_n31), .S(
        MULi_5_mult_15_n28), .ICO(MULi_5_mult_15_n26), .CO(MULi_5_mult_15_n27)
         );
  CMPR42X1 MULi_5_mult_15_U20 ( .A(MULi_5_mult_15_n72), .B(MULi_5_mult_15_n65), 
        .C(MULi_5_mult_15_n59), .D(n162), .ICI(MULi_5_mult_15_n26), .S(
        MULi_5_mult_15_n25), .ICO(MULi_5_mult_15_n23), .CO(MULi_5_mult_15_n24)
         );
  ADDFX1 MULi_6_mult_15_U5 ( .A(MULi_6_mult_15_n24), .B(MULi_6_mult_15_n20), 
        .CI(MULi_6_mult_15_n5), .CO(MULi_6_mult_15_n4), .S(MUL_to_PIPE1[11])
         );
  ADDFX1 MULi_6_mult_15_U6 ( .A(MULi_6_mult_15_n27), .B(MULi_6_mult_15_n25), 
        .CI(MULi_6_mult_15_n6), .CO(MULi_6_mult_15_n5), .S(MUL_to_PIPE1[10])
         );
  ADDFX1 MULi_6_mult_15_U7 ( .A(MULi_6_mult_15_n28), .B(MULi_6_mult_15_n32), 
        .CI(MULi_6_mult_15_n7), .CO(MULi_6_mult_15_n6), .S(MUL_to_PIPE1[9]) );
  ADDFX1 MULi_6_mult_15_U8 ( .A(MULi_6_mult_15_n33), .B(MULi_6_mult_15_n37), 
        .CI(MULi_6_mult_15_n8), .CO(MULi_6_mult_15_n7), .S(MUL_to_PIPE1[8]) );
  ADDFX1 MULi_6_mult_15_U9 ( .A(MULi_6_mult_15_n38), .B(MULi_6_mult_15_n42), 
        .CI(MULi_6_mult_15_n9), .CO(MULi_6_mult_15_n8), .S(MUL_to_PIPE1[7]) );
  ADDFX1 MULi_6_mult_15_U10 ( .A(MULi_6_mult_15_n44), .B(MULi_6_mult_15_n43), 
        .CI(MULi_6_mult_15_n10), .CO(MULi_6_mult_15_n9), .S(MUL_to_PIPE1[6])
         );
  ADDFX1 MULi_6_mult_15_U11 ( .A(MULi_6_mult_15_n45), .B(MULi_6_mult_15_n47), 
        .CI(MULi_6_mult_15_n11), .CO(MULi_6_mult_15_n10), .S(MUL_to_PIPE1[5])
         );
  ADDFX1 MULi_6_mult_15_U12 ( .A(MULi_6_mult_15_n49), .B(MULi_6_mult_15_n50), 
        .CI(MULi_6_mult_15_n12), .CO(MULi_6_mult_15_n11), .S(MUL_to_PIPE1[4])
         );
  ADDFX1 MULi_6_mult_15_U13 ( .A(MULi_6_mult_15_n51), .B(MULi_6_mult_15_n54), 
        .CI(MULi_6_mult_15_n13), .CO(MULi_6_mult_15_n12), .S(MUL_to_PIPE1[3])
         );
  ADDFX1 MULi_6_mult_15_U14 ( .A(MULi_6_mult_15_n86), .B(MULi_6_mult_15_n79), 
        .CI(MULi_6_mult_15_n14), .CO(MULi_6_mult_15_n13), .S(MUL_to_PIPE1[2])
         );
  ADDHX1 MULi_6_mult_15_U15 ( .A(MULi_6_mult_15_n55), .B(MULi_6_mult_15_n87), 
        .CO(MULi_6_mult_15_n14), .S(MUL_to_PIPE1[1]) );
  ADDFX1 MULi_6_mult_15_U29 ( .A(MULi_6_mult_15_n70), .B(MULi_6_mult_15_n76), 
        .CI(MULi_6_mult_15_n48), .CO(MULi_6_mult_15_n44), .S(
        MULi_6_mult_15_n45) );
  ADDFX1 MULi_6_mult_15_U31 ( .A(MULi_6_mult_15_n84), .B(MULi_6_mult_15_n71), 
        .CI(MULi_6_mult_15_n77), .CO(MULi_6_mult_15_n48), .S(
        MULi_6_mult_15_n49) );
  ADDFX1 MULi_6_mult_15_U18 ( .A(MULi_6_mult_15_n22), .B(MULi_6_mult_15_n58), 
        .CI(MULi_6_mult_15_n23), .CO(MULi_6_mult_15_n19), .S(
        MULi_6_mult_15_n20) );
  ADDFX1 MULi_6_mult_15_U17 ( .A(MULi_6_mult_15_n57), .B(MULi_6_mult_15_n64), 
        .CI(MULi_6_mult_15_n21), .CO(MULi_6_mult_15_n17), .S(
        MULi_6_mult_15_n18) );
  CMPR42X1 MULi_6_mult_15_U28 ( .A(MULi_6_mult_15_n63), .B(MULi_6_mult_15_n82), 
        .C(MULi_6_mult_15_n75), .D(MULi_6_mult_15_n69), .ICI(
        MULi_6_mult_15_n46), .S(MULi_6_mult_15_n43), .ICO(MULi_6_mult_15_n41), 
        .CO(MULi_6_mult_15_n42) );
  CMPR42X1 MULi_6_mult_15_U26 ( .A(MULi_6_mult_15_n74), .B(MULi_6_mult_15_n62), 
        .C(MULi_6_mult_15_n68), .D(MULi_6_mult_15_n41), .ICI(
        MULi_6_mult_15_n40), .S(MULi_6_mult_15_n38), .ICO(MULi_6_mult_15_n36), 
        .CO(MULi_6_mult_15_n37) );
  CMPR42X1 MULi_6_mult_15_U23 ( .A(MULi_6_mult_15_n67), .B(MULi_6_mult_15_n61), 
        .C(MULi_6_mult_15_n39), .D(MULi_6_mult_15_n36), .ICI(
        MULi_6_mult_15_n35), .S(MULi_6_mult_15_n33), .ICO(MULi_6_mult_15_n31), 
        .CO(MULi_6_mult_15_n32) );
  CMPR42X1 MULi_6_mult_15_U21 ( .A(MULi_6_mult_15_n66), .B(MULi_6_mult_15_n60), 
        .C(n157), .D(MULi_6_mult_15_n34), .ICI(MULi_6_mult_15_n31), .S(
        MULi_6_mult_15_n28), .ICO(MULi_6_mult_15_n26), .CO(MULi_6_mult_15_n27)
         );
  CMPR42X1 MULi_6_mult_15_U20 ( .A(MULi_6_mult_15_n72), .B(MULi_6_mult_15_n65), 
        .C(MULi_6_mult_15_n59), .D(n156), .ICI(MULi_6_mult_15_n26), .S(
        MULi_6_mult_15_n25), .ICO(MULi_6_mult_15_n23), .CO(MULi_6_mult_15_n24)
         );
  ADDFX1 MULi_0_mult_15_U2 ( .A(MULi_0_mult_15_n15), .B(MULi_0_mult_15_n56), 
        .CI(MULi_0_mult_15_n2), .CO(MULi_0_mult_15_n1), .S(MUL_to_PIPE1[110])
         );
  ADDFX1 MULi_0_mult_15_U3 ( .A(MULi_0_mult_15_n17), .B(MULi_0_mult_15_n16), 
        .CI(MULi_0_mult_15_n3), .CO(MULi_0_mult_15_n2), .S(MUL_to_PIPE1[109])
         );
  ADDFX1 MULi_0_mult_15_U4 ( .A(MULi_0_mult_15_n19), .B(MULi_0_mult_15_n18), 
        .CI(MULi_0_mult_15_n4), .CO(MULi_0_mult_15_n3), .S(MUL_to_PIPE1[108])
         );
  ADDFX1 MULi_0_mult_15_U5 ( .A(MULi_0_mult_15_n24), .B(MULi_0_mult_15_n20), 
        .CI(MULi_0_mult_15_n5), .CO(MULi_0_mult_15_n4), .S(MUL_to_PIPE1[107])
         );
  ADDFX1 MULi_0_mult_15_U6 ( .A(MULi_0_mult_15_n27), .B(MULi_0_mult_15_n25), 
        .CI(MULi_0_mult_15_n6), .CO(MULi_0_mult_15_n5), .S(MUL_to_PIPE1[106])
         );
  ADDFX1 MULi_0_mult_15_U7 ( .A(MULi_0_mult_15_n28), .B(MULi_0_mult_15_n32), 
        .CI(MULi_0_mult_15_n7), .CO(MULi_0_mult_15_n6), .S(MUL_to_PIPE1[105])
         );
  ADDFX1 MULi_0_mult_15_U8 ( .A(MULi_0_mult_15_n33), .B(MULi_0_mult_15_n37), 
        .CI(MULi_0_mult_15_n8), .CO(MULi_0_mult_15_n7), .S(MUL_to_PIPE1[104])
         );
  ADDFX1 MULi_0_mult_15_U9 ( .A(MULi_0_mult_15_n38), .B(MULi_0_mult_15_n42), 
        .CI(MULi_0_mult_15_n9), .CO(MULi_0_mult_15_n8), .S(MUL_to_PIPE1[103])
         );
  ADDFX1 MULi_0_mult_15_U10 ( .A(MULi_0_mult_15_n44), .B(MULi_0_mult_15_n43), 
        .CI(MULi_0_mult_15_n10), .CO(MULi_0_mult_15_n9), .S(MUL_to_PIPE1[102])
         );
  ADDFX1 MULi_0_mult_15_U11 ( .A(MULi_0_mult_15_n45), .B(MULi_0_mult_15_n47), 
        .CI(MULi_0_mult_15_n11), .CO(MULi_0_mult_15_n10), .S(MUL_to_PIPE1[101]) );
  ADDFX1 MULi_0_mult_15_U12 ( .A(MULi_0_mult_15_n49), .B(MULi_0_mult_15_n50), 
        .CI(MULi_0_mult_15_n12), .CO(MULi_0_mult_15_n11), .S(MUL_to_PIPE1[100]) );
  ADDFX1 MULi_0_mult_15_U13 ( .A(MULi_0_mult_15_n51), .B(MULi_0_mult_15_n54), 
        .CI(MULi_0_mult_15_n13), .CO(MULi_0_mult_15_n12), .S(MUL_to_PIPE1[99])
         );
  ADDFX1 MULi_0_mult_15_U14 ( .A(MULi_0_mult_15_n86), .B(MULi_0_mult_15_n79), 
        .CI(MULi_0_mult_15_n14), .CO(MULi_0_mult_15_n13), .S(MUL_to_PIPE1[98])
         );
  ADDHX1 MULi_0_mult_15_U15 ( .A(MULi_0_mult_15_n55), .B(MULi_0_mult_15_n87), 
        .CO(MULi_0_mult_15_n14), .S(MUL_to_PIPE1[97]) );
  ADDFX1 MULi_0_mult_15_U29 ( .A(MULi_0_mult_15_n70), .B(MULi_0_mult_15_n76), 
        .CI(MULi_0_mult_15_n48), .CO(MULi_0_mult_15_n44), .S(
        MULi_0_mult_15_n45) );
  ADDFX1 MULi_0_mult_15_U31 ( .A(MULi_0_mult_15_n84), .B(MULi_0_mult_15_n71), 
        .CI(MULi_0_mult_15_n77), .CO(MULi_0_mult_15_n48), .S(
        MULi_0_mult_15_n49) );
  ADDFX1 MULi_0_mult_15_U18 ( .A(MULi_0_mult_15_n22), .B(MULi_0_mult_15_n58), 
        .CI(MULi_0_mult_15_n23), .CO(MULi_0_mult_15_n19), .S(
        MULi_0_mult_15_n20) );
  ADDFX1 MULi_0_mult_15_U17 ( .A(MULi_0_mult_15_n57), .B(MULi_0_mult_15_n64), 
        .CI(MULi_0_mult_15_n21), .CO(MULi_0_mult_15_n17), .S(
        MULi_0_mult_15_n18) );
  CMPR42X1 MULi_0_mult_15_U28 ( .A(MULi_0_mult_15_n63), .B(MULi_0_mult_15_n82), 
        .C(MULi_0_mult_15_n75), .D(MULi_0_mult_15_n69), .ICI(
        MULi_0_mult_15_n46), .S(MULi_0_mult_15_n43), .ICO(MULi_0_mult_15_n41), 
        .CO(MULi_0_mult_15_n42) );
  CMPR42X1 MULi_0_mult_15_U26 ( .A(MULi_0_mult_15_n74), .B(MULi_0_mult_15_n62), 
        .C(MULi_0_mult_15_n68), .D(MULi_0_mult_15_n41), .ICI(
        MULi_0_mult_15_n40), .S(MULi_0_mult_15_n38), .ICO(MULi_0_mult_15_n36), 
        .CO(MULi_0_mult_15_n37) );
  CMPR42X1 MULi_0_mult_15_U23 ( .A(MULi_0_mult_15_n67), .B(MULi_0_mult_15_n61), 
        .C(MULi_0_mult_15_n39), .D(MULi_0_mult_15_n36), .ICI(
        MULi_0_mult_15_n35), .S(MULi_0_mult_15_n33), .ICO(MULi_0_mult_15_n31), 
        .CO(MULi_0_mult_15_n32) );
  CMPR42X1 MULi_0_mult_15_U21 ( .A(MULi_0_mult_15_n66), .B(MULi_0_mult_15_n60), 
        .C(n167), .D(MULi_0_mult_15_n34), .ICI(MULi_0_mult_15_n31), .S(
        MULi_0_mult_15_n28), .ICO(MULi_0_mult_15_n26), .CO(MULi_0_mult_15_n27)
         );
  CMPR42X1 MULi_0_mult_15_U20 ( .A(MULi_0_mult_15_n72), .B(MULi_0_mult_15_n65), 
        .C(MULi_0_mult_15_n59), .D(n166), .ICI(MULi_0_mult_15_n26), .S(
        MULi_0_mult_15_n25), .ICO(MULi_0_mult_15_n23), .CO(MULi_0_mult_15_n24)
         );
  AND2X2 U66 ( .A(VIN), .B(SR_to_MUX), .Y(MUX_to_PIPE1) );
  OR2X2 U57 ( .A(VIN), .B(SR_SRI_bit_temp_out[0]), .Y(n62) );
  DFFRX4 REG_IN_H_i_6_q_reg_7_ ( .D(H6[7]), .CK(CLK), .RN(RST_n), .Q(TEMP_H[7]), .QN(n336) );
  DFFRX4 REG_IN_H_i_6_q_reg_6_ ( .D(H6[6]), .CK(CLK), .RN(RST_n), .Q(TEMP_H[6]), .QN(n338) );
  DFFRX4 REG_IN_H_i_6_q_reg_5_ ( .D(H6[5]), .CK(CLK), .RN(RST_n), .Q(TEMP_H[5]), .QN(n340) );
  DFFRX4 REG_IN_H_i_6_q_reg_4_ ( .D(H6[4]), .CK(CLK), .RN(RST_n), .Q(TEMP_H[4]), .QN(n342) );
  DFFRX4 REG_IN_H_i_6_q_reg_3_ ( .D(H6[3]), .CK(CLK), .RN(RST_n), .Q(TEMP_H[3]), .QN(n344) );
  DFFRX4 REG_IN_H_i_6_q_reg_2_ ( .D(H6[2]), .CK(CLK), .RN(RST_n), .Q(TEMP_H[2]), .QN(n346) );
  DFFRX4 REG_IN_H_i_6_q_reg_0_ ( .D(H6[0]), .CK(CLK), .RN(RST_n), .Q(TEMP_H[0]), .QN(n351) );
  DFFRX4 REG_IN_H_i_5_q_reg_7_ ( .D(H5[7]), .CK(CLK), .RN(RST_n), .Q(
        TEMP_H[15]), .QN(n400) );
  DFFRX4 REG_IN_H_i_5_q_reg_6_ ( .D(H5[6]), .CK(CLK), .RN(RST_n), .Q(
        TEMP_H[14]), .QN(n402) );
  DFFRX4 REG_IN_H_i_5_q_reg_5_ ( .D(H5[5]), .CK(CLK), .RN(RST_n), .Q(
        TEMP_H[13]), .QN(n404) );
  DFFRX4 REG_IN_H_i_5_q_reg_4_ ( .D(H5[4]), .CK(CLK), .RN(RST_n), .Q(
        TEMP_H[12]), .QN(n406) );
  DFFRX4 REG_IN_H_i_5_q_reg_3_ ( .D(H5[3]), .CK(CLK), .RN(RST_n), .Q(
        TEMP_H[11]), .QN(n408) );
  DFFRX4 REG_IN_H_i_5_q_reg_2_ ( .D(H5[2]), .CK(CLK), .RN(RST_n), .Q(
        TEMP_H[10]), .QN(n410) );
  DFFRX4 REG_IN_H_i_5_q_reg_0_ ( .D(H5[0]), .CK(CLK), .RN(RST_n), .Q(TEMP_H[8]), .QN(n415) );
  DFFRX4 REG_IN_H_i_4_q_reg_7_ ( .D(H4[7]), .CK(CLK), .RN(RST_n), .Q(
        TEMP_H[23]), .QN(n464) );
  DFFRX4 REG_IN_H_i_4_q_reg_6_ ( .D(H4[6]), .CK(CLK), .RN(RST_n), .Q(
        TEMP_H[22]), .QN(n466) );
  DFFRX4 REG_IN_H_i_4_q_reg_5_ ( .D(H4[5]), .CK(CLK), .RN(RST_n), .Q(
        TEMP_H[21]), .QN(n468) );
  DFFRX4 REG_IN_H_i_4_q_reg_4_ ( .D(H4[4]), .CK(CLK), .RN(RST_n), .Q(
        TEMP_H[20]), .QN(n470) );
  DFFRX4 REG_IN_H_i_4_q_reg_3_ ( .D(H4[3]), .CK(CLK), .RN(RST_n), .Q(
        TEMP_H[19]), .QN(n472) );
  DFFRX4 REG_IN_H_i_4_q_reg_2_ ( .D(H4[2]), .CK(CLK), .RN(RST_n), .Q(
        TEMP_H[18]), .QN(n474) );
  DFFRX4 REG_IN_H_i_4_q_reg_0_ ( .D(H4[0]), .CK(CLK), .RN(RST_n), .Q(
        TEMP_H[16]), .QN(n479) );
  DFFRX4 REG_IN_H_i_3_q_reg_7_ ( .D(H3[7]), .CK(CLK), .RN(RST_n), .Q(
        TEMP_H[31]), .QN(n528) );
  DFFRX4 REG_IN_H_i_3_q_reg_6_ ( .D(H3[6]), .CK(CLK), .RN(RST_n), .Q(
        TEMP_H[30]), .QN(n530) );
  DFFRX4 REG_IN_H_i_3_q_reg_5_ ( .D(H3[5]), .CK(CLK), .RN(RST_n), .Q(
        TEMP_H[29]), .QN(n532) );
  DFFRX4 REG_IN_H_i_3_q_reg_4_ ( .D(H3[4]), .CK(CLK), .RN(RST_n), .Q(
        TEMP_H[28]), .QN(n534) );
  DFFRX4 REG_IN_H_i_3_q_reg_3_ ( .D(H3[3]), .CK(CLK), .RN(RST_n), .Q(
        TEMP_H[27]), .QN(n536) );
  DFFRX4 REG_IN_H_i_3_q_reg_2_ ( .D(H3[2]), .CK(CLK), .RN(RST_n), .Q(
        TEMP_H[26]), .QN(n538) );
  DFFRX4 REG_IN_H_i_3_q_reg_0_ ( .D(H3[0]), .CK(CLK), .RN(RST_n), .Q(
        TEMP_H[24]), .QN(n543) );
  DFFRX4 REG_IN_H_i_2_q_reg_7_ ( .D(H2[7]), .CK(CLK), .RN(RST_n), .Q(
        TEMP_H[39]), .QN(n592) );
  DFFRX4 REG_IN_H_i_2_q_reg_6_ ( .D(H2[6]), .CK(CLK), .RN(RST_n), .Q(
        TEMP_H[38]), .QN(n594) );
  DFFRX4 REG_IN_H_i_2_q_reg_5_ ( .D(H2[5]), .CK(CLK), .RN(RST_n), .Q(
        TEMP_H[37]), .QN(n596) );
  DFFRX4 REG_IN_H_i_2_q_reg_4_ ( .D(H2[4]), .CK(CLK), .RN(RST_n), .Q(
        TEMP_H[36]), .QN(n598) );
  DFFRX4 REG_IN_H_i_2_q_reg_3_ ( .D(H2[3]), .CK(CLK), .RN(RST_n), .Q(
        TEMP_H[35]), .QN(n600) );
  DFFRX4 REG_IN_H_i_2_q_reg_2_ ( .D(H2[2]), .CK(CLK), .RN(RST_n), .Q(
        TEMP_H[34]), .QN(n602) );
  DFFRX4 REG_IN_H_i_2_q_reg_0_ ( .D(H2[0]), .CK(CLK), .RN(RST_n), .Q(
        TEMP_H[32]), .QN(n607) );
  DFFRX4 REG_IN_H_i_1_q_reg_7_ ( .D(H1[7]), .CK(CLK), .RN(RST_n), .Q(
        TEMP_H[47]), .QN(n656) );
  DFFRX4 REG_IN_H_i_1_q_reg_6_ ( .D(H1[6]), .CK(CLK), .RN(RST_n), .Q(
        TEMP_H[46]), .QN(n658) );
  DFFRX4 REG_IN_H_i_1_q_reg_5_ ( .D(H1[5]), .CK(CLK), .RN(RST_n), .Q(
        TEMP_H[45]), .QN(n660) );
  DFFRX4 REG_IN_H_i_1_q_reg_4_ ( .D(H1[4]), .CK(CLK), .RN(RST_n), .Q(
        TEMP_H[44]), .QN(n662) );
  DFFRX4 REG_IN_H_i_1_q_reg_3_ ( .D(H1[3]), .CK(CLK), .RN(RST_n), .Q(
        TEMP_H[43]), .QN(n664) );
  DFFRX4 REG_IN_H_i_1_q_reg_2_ ( .D(H1[2]), .CK(CLK), .RN(RST_n), .Q(
        TEMP_H[42]), .QN(n666) );
  DFFRX4 REG_IN_H_i_1_q_reg_0_ ( .D(H1[0]), .CK(CLK), .RN(RST_n), .Q(
        TEMP_H[40]), .QN(n671) );
  DFFRX4 REG_IN_H_i_0_q_reg_7_ ( .D(H0[7]), .CK(CLK), .RN(RST_n), .Q(
        TEMP_H[55]), .QN(n272) );
  DFFRX4 REG_IN_H_i_0_q_reg_6_ ( .D(H0[6]), .CK(CLK), .RN(RST_n), .Q(
        TEMP_H[54]), .QN(n274) );
  DFFRX4 REG_IN_H_i_0_q_reg_5_ ( .D(H0[5]), .CK(CLK), .RN(RST_n), .Q(
        TEMP_H[53]), .QN(n276) );
  DFFRX4 REG_IN_H_i_0_q_reg_4_ ( .D(H0[4]), .CK(CLK), .RN(RST_n), .Q(
        TEMP_H[52]), .QN(n278) );
  DFFRX4 REG_IN_H_i_0_q_reg_3_ ( .D(H0[3]), .CK(CLK), .RN(RST_n), .Q(
        TEMP_H[51]), .QN(n280) );
  DFFRX4 REG_IN_H_i_0_q_reg_2_ ( .D(H0[2]), .CK(CLK), .RN(RST_n), .Q(
        TEMP_H[50]), .QN(n282) );
  DFFRX4 REG_IN_H_i_0_q_reg_0_ ( .D(H0[0]), .CK(CLK), .RN(RST_n), .Q(
        TEMP_H[48]), .QN(n287) );
  DFFRX4 REG_IN_H_i_6_q_reg_1_ ( .D(H6[1]), .CK(CLK), .RN(RST_n), .Q(TEMP_H[1]), .QN(n347) );
  DFFRX4 REG_IN_H_i_5_q_reg_1_ ( .D(H5[1]), .CK(CLK), .RN(RST_n), .Q(TEMP_H[9]), .QN(n411) );
  DFFRX4 REG_IN_H_i_4_q_reg_1_ ( .D(H4[1]), .CK(CLK), .RN(RST_n), .Q(
        TEMP_H[17]), .QN(n475) );
  DFFRX4 REG_IN_H_i_3_q_reg_1_ ( .D(H3[1]), .CK(CLK), .RN(RST_n), .Q(
        TEMP_H[25]), .QN(n539) );
  DFFRX4 REG_IN_H_i_2_q_reg_1_ ( .D(H2[1]), .CK(CLK), .RN(RST_n), .Q(
        TEMP_H[33]), .QN(n603) );
  DFFRX4 REG_IN_H_i_1_q_reg_1_ ( .D(H1[1]), .CK(CLK), .RN(RST_n), .Q(
        TEMP_H[41]), .QN(n667) );
  DFFRX4 REG_IN_H_i_0_q_reg_1_ ( .D(H0[1]), .CK(CLK), .RN(RST_n), .Q(
        TEMP_H[49]), .QN(n283) );
  DFFRX4 SR_SRI_regi_6_q_reg_0_ ( .D(n50), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[0]), .QN(n352) );
  DFFRX4 SR_SRI_regi_5_q_reg_0_ ( .D(n51), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[8]), .QN(n416) );
  DFFRX4 SR_SRI_regi_4_q_reg_0_ ( .D(n52), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[16]), .QN(n480) );
  DFFRX4 SR_SRI_regi_3_q_reg_0_ ( .D(n53), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[24]), .QN(n544) );
  DFFRX4 SR_SRI_regi_2_q_reg_0_ ( .D(n54), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[32]), .QN(n608) );
  DFFRX4 SR_SRI_regi_1_q_reg_0_ ( .D(n55), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[40]), .QN(n672) );
  DFFRX4 SR_SRI_reg0_q_reg_0_ ( .D(n70), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[48]), .QN(n288) );
  DFFRX4 SR_SRI_regi_5_q_reg_7_ ( .D(n9), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[15]) );
  DFFRX4 SR_SRI_regi_5_q_reg_5_ ( .D(n21), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[13]) );
  DFFRX4 SR_SRI_regi_5_q_reg_3_ ( .D(n33), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[11]) );
  DFFRX4 SR_SRI_regi_5_q_reg_1_ ( .D(n45), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[9]) );
  DFFRX4 SR_SRI_regi_4_q_reg_7_ ( .D(n10), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[23]) );
  DFFRX4 SR_SRI_regi_4_q_reg_5_ ( .D(n22), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[21]) );
  DFFRX4 SR_SRI_regi_4_q_reg_3_ ( .D(n34), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[19]) );
  DFFRX4 SR_SRI_regi_4_q_reg_1_ ( .D(n46), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[17]) );
  DFFRX4 SR_SRI_regi_3_q_reg_7_ ( .D(n11), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[31]) );
  DFFRX4 SR_SRI_regi_3_q_reg_5_ ( .D(n23), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[29]) );
  DFFRX4 SR_SRI_regi_3_q_reg_3_ ( .D(n35), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[27]) );
  DFFRX4 SR_SRI_regi_3_q_reg_1_ ( .D(n47), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[25]) );
  DFFRX4 SR_SRI_regi_2_q_reg_7_ ( .D(n12), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[39]) );
  DFFRX4 SR_SRI_regi_2_q_reg_5_ ( .D(n24), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[37]) );
  DFFRX4 SR_SRI_regi_2_q_reg_3_ ( .D(n36), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[35]) );
  DFFRX4 SR_SRI_regi_2_q_reg_1_ ( .D(n48), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[33]) );
  DFFRX4 SR_SRI_regi_1_q_reg_7_ ( .D(n13), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[47]) );
  DFFRX4 SR_SRI_regi_1_q_reg_5_ ( .D(n25), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[45]) );
  DFFRX4 SR_SRI_regi_1_q_reg_3_ ( .D(n37), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[43]) );
  DFFRX4 SR_SRI_regi_1_q_reg_1_ ( .D(n49), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[41]) );
  DFFRX4 SR_SRI_reg0_q_reg_7_ ( .D(n63), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[55]) );
  DFFRX4 SR_SRI_reg0_q_reg_5_ ( .D(n65), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[53]) );
  DFFRX4 SR_SRI_reg0_q_reg_3_ ( .D(n67), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[51]) );
  DFFRX4 SR_SRI_reg0_q_reg_1_ ( .D(n69), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[49]) );
  DFFRX4 SR_SRI_regi_6_q_reg_6_ ( .D(n14), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[6]), .QN(n297) );
  DFFRX4 SR_SRI_regi_6_q_reg_4_ ( .D(n26), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[4]), .QN(n298) );
  DFFRX4 SR_SRI_regi_5_q_reg_6_ ( .D(n15), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[14]), .QN(n361) );
  DFFRX4 SR_SRI_regi_5_q_reg_4_ ( .D(n27), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[12]), .QN(n362) );
  DFFRX4 SR_SRI_regi_5_q_reg_2_ ( .D(n39), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[10]), .QN(n363) );
  DFFRX4 SR_SRI_regi_4_q_reg_6_ ( .D(n16), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[22]), .QN(n425) );
  DFFRX4 SR_SRI_regi_4_q_reg_4_ ( .D(n28), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[20]), .QN(n426) );
  DFFRX4 SR_SRI_regi_4_q_reg_2_ ( .D(n40), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[18]), .QN(n427) );
  DFFRX4 SR_SRI_regi_3_q_reg_6_ ( .D(n17), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[30]), .QN(n489) );
  DFFRX4 SR_SRI_regi_3_q_reg_4_ ( .D(n29), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[28]), .QN(n490) );
  DFFRX4 SR_SRI_regi_3_q_reg_2_ ( .D(n41), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[26]), .QN(n491) );
  DFFRX4 SR_SRI_regi_2_q_reg_6_ ( .D(n18), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[38]), .QN(n553) );
  DFFRX4 SR_SRI_regi_2_q_reg_4_ ( .D(n30), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[36]), .QN(n554) );
  DFFRX4 SR_SRI_regi_2_q_reg_2_ ( .D(n42), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[34]), .QN(n555) );
  DFFRX4 SR_SRI_regi_1_q_reg_6_ ( .D(n19), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[46]), .QN(n617) );
  DFFRX4 SR_SRI_regi_1_q_reg_4_ ( .D(n31), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[44]), .QN(n618) );
  DFFRX4 SR_SRI_regi_1_q_reg_2_ ( .D(n43), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[42]), .QN(n619) );
  DFFRX4 SR_SRI_reg0_q_reg_6_ ( .D(n64), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[54]), .QN(n233) );
  DFFRX4 SR_SRI_reg0_q_reg_4_ ( .D(n66), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[52]), .QN(n234) );
  DFFRX4 SR_SRI_reg0_q_reg_2_ ( .D(n68), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[50]), .QN(n235) );
  DFFRX4 SR_SRI_regi_6_q_reg_2_ ( .D(n38), .CK(CLK), .RN(RST_n), .Q(
        SR_to_MUL[2]), .QN(n299) );
  OAI2BB2X4 U67 ( .B0(n73), .B1(n687), .A0N(ADD_esteso_13__7_), .A1N(
        ADD_esteso_12__7_), .Y(n688) );
  OAI2BB2X4 U68 ( .B0(n72), .B1(n685), .A0N(ADD_esteso_13__5_), .A1N(
        ADD_esteso_12__5_), .Y(n686) );
  OAI2BB2X4 U69 ( .B0(n71), .B1(n683), .A0N(ADD_esteso_13__3_), .A1N(
        ADD_esteso_12__3_), .Y(n684) );
  OR2X8 U70 ( .A(n227), .B(n228), .Y(n75) );
  OR2X8 U71 ( .A(n221), .B(n222), .Y(n78) );
  OR2X8 U72 ( .A(n223), .B(n224), .Y(n77) );
  OR2X8 U73 ( .A(n219), .B(n220), .Y(n79) );
  OR2X8 U74 ( .A(n225), .B(n226), .Y(n76) );
  OR2X8 U75 ( .A(n231), .B(n232), .Y(n80) );
  OR2X8 U76 ( .A(n229), .B(n230), .Y(n74) );
  NOR2X2 U77 ( .A(ADD_esteso_13__3_), .B(ADD_esteso_12__3_), .Y(n71) );
  NOR2X2 U78 ( .A(ADD_esteso_13__5_), .B(ADD_esteso_12__5_), .Y(n72) );
  NOR2X2 U79 ( .A(ADD_esteso_13__7_), .B(ADD_esteso_12__7_), .Y(n73) );
  NAND2X2 U80 ( .A(n676), .B(n672), .Y(n670) );
  NAND2X2 U81 ( .A(n612), .B(n608), .Y(n606) );
  NAND2X2 U82 ( .A(n420), .B(n416), .Y(n414) );
  CLKNAND2X2 U83 ( .A(n356), .B(n352), .Y(n350) );
  NAND2X2 U84 ( .A(n292), .B(n288), .Y(n286) );
  NAND2X2 U85 ( .A(n548), .B(n544), .Y(n542) );
  NAND2X2 U86 ( .A(n484), .B(n480), .Y(n478) );
  INVX16 U87 ( .A(n354), .Y(n320) );
  AOI22X1 U88 ( .A0(n356), .A1(n338), .B0(n93), .B1(n150), .Y(n339) );
  AOI22X1 U89 ( .A0(n95), .A1(n309), .B0(n353), .B1(n342), .Y(n306) );
  OAI22X1 U90 ( .A0(n359), .A1(n316), .B0(n360), .B1(n317), .Y(
        MULi_6_mult_15_n66) );
  ADDHX2 U91 ( .A(MULi_4_mult_15_n85), .B(MULi_4_mult_15_n78), .CO(
        MULi_4_mult_15_n50), .S(MULi_4_mult_15_n51) );
  OAI22X1 U92 ( .A0(n78), .A1(n463), .B0(n462), .B1(n461), .Y(
        MULi_4_mult_15_n78) );
  ADDHX2 U93 ( .A(MULi_5_mult_15_n85), .B(MULi_5_mult_15_n78), .CO(
        MULi_5_mult_15_n50), .S(MULi_5_mult_15_n51) );
  OAI22X1 U94 ( .A0(n79), .A1(n399), .B0(n398), .B1(n397), .Y(
        MULi_5_mult_15_n78) );
  ADDHX2 U95 ( .A(MULi_2_mult_15_n85), .B(MULi_2_mult_15_n78), .CO(
        MULi_2_mult_15_n50), .S(MULi_2_mult_15_n51) );
  OAI22X1 U96 ( .A0(n77), .A1(n591), .B0(n590), .B1(n589), .Y(
        MULi_2_mult_15_n78) );
  ADDHX2 U97 ( .A(MULi_0_mult_15_n85), .B(MULi_0_mult_15_n78), .CO(
        MULi_0_mult_15_n50), .S(MULi_0_mult_15_n51) );
  OAI22X1 U98 ( .A0(n76), .A1(n271), .B0(n270), .B1(n269), .Y(
        MULi_0_mult_15_n78) );
  ADDHX2 U99 ( .A(MULi_3_mult_15_n85), .B(MULi_3_mult_15_n78), .CO(
        MULi_3_mult_15_n50), .S(MULi_3_mult_15_n51) );
  OAI22X1 U100 ( .A0(n74), .A1(n527), .B0(n526), .B1(n525), .Y(
        MULi_3_mult_15_n78) );
  ADDHX2 U101 ( .A(MULi_6_mult_15_n85), .B(MULi_6_mult_15_n78), .CO(
        MULi_6_mult_15_n50), .S(MULi_6_mult_15_n51) );
  OAI22X1 U102 ( .A0(n80), .A1(n335), .B0(n334), .B1(n333), .Y(
        MULi_6_mult_15_n78) );
  ADDHX2 U103 ( .A(MULi_1_mult_15_n85), .B(MULi_1_mult_15_n78), .CO(
        MULi_1_mult_15_n50), .S(MULi_1_mult_15_n51) );
  AOI22X1 U104 ( .A0(n548), .A1(n534), .B0(TEMP_H[28]), .B1(n152), .Y(n535) );
  AOI22X1 U105 ( .A0(n548), .A1(n536), .B0(TEMP_H[27]), .B1(n152), .Y(n537) );
  AOI22X1 U106 ( .A0(n612), .A1(n600), .B0(TEMP_H[35]), .B1(n153), .Y(n601) );
  AOI22X1 U107 ( .A0(n484), .A1(n470), .B0(TEMP_H[20]), .B1(n154), .Y(n471) );
  AOI22X1 U108 ( .A0(n612), .A1(n598), .B0(TEMP_H[36]), .B1(n153), .Y(n599) );
  AOI22X1 U109 ( .A0(n484), .A1(n472), .B0(TEMP_H[19]), .B1(n154), .Y(n473) );
  AOI22X1 U110 ( .A0(n676), .A1(n664), .B0(TEMP_H[43]), .B1(n148), .Y(n665) );
  AOI22X1 U111 ( .A0(n420), .A1(n406), .B0(TEMP_H[12]), .B1(n151), .Y(n407) );
  AOI22X1 U112 ( .A0(n676), .A1(n662), .B0(TEMP_H[44]), .B1(n148), .Y(n663) );
  AOI22X1 U113 ( .A0(n420), .A1(n408), .B0(TEMP_H[11]), .B1(n151), .Y(n409) );
  AOI22X1 U114 ( .A0(n292), .A1(n280), .B0(TEMP_H[51]), .B1(n149), .Y(n281) );
  AOI22X1 U115 ( .A0(n356), .A1(n344), .B0(TEMP_H[3]), .B1(n150), .Y(n345) );
  AOI22X1 U116 ( .A0(n292), .A1(n278), .B0(TEMP_H[52]), .B1(n149), .Y(n279) );
  CLKINVX2 U117 ( .A(n532), .Y(n81) );
  CLKINVX2 U118 ( .A(n596), .Y(n82) );
  CLKINVX2 U119 ( .A(n468), .Y(n83) );
  CLKINVX2 U120 ( .A(n660), .Y(n84) );
  CLKINVX2 U121 ( .A(n404), .Y(n85) );
  CLKINVX2 U122 ( .A(n276), .Y(n86) );
  CLKINVX2 U123 ( .A(n340), .Y(n87) );
  INVX1 U124 ( .A(n530), .Y(n88) );
  INVX1 U125 ( .A(n466), .Y(n89) );
  INVX1 U126 ( .A(n594), .Y(n90) );
  INVX1 U127 ( .A(n402), .Y(n91) );
  INVX1 U128 ( .A(n658), .Y(n92) );
  INVX1 U129 ( .A(n338), .Y(n93) );
  INVX1 U130 ( .A(n274), .Y(n94) );
  BUFX2 U131 ( .A(TEMP_H[4]), .Y(n95) );
  CLKINVX2 U132 ( .A(n105), .Y(n96) );
  CLKBUFX6 U133 ( .A(TEMP_H[16]), .Y(n105) );
  CLKINVX2 U134 ( .A(n107), .Y(n97) );
  CLKBUFX6 U135 ( .A(TEMP_H[8]), .Y(n107) );
  CLKINVX2 U136 ( .A(n104), .Y(n98) );
  CLKBUFX6 U137 ( .A(TEMP_H[24]), .Y(n104) );
  CLKINVX2 U138 ( .A(n109), .Y(n99) );
  CLKBUFX6 U139 ( .A(TEMP_H[0]), .Y(n109) );
  CLKINVX2 U140 ( .A(n106), .Y(n100) );
  CLKBUFX6 U141 ( .A(TEMP_H[32]), .Y(n106) );
  CLKINVX2 U142 ( .A(n110), .Y(n101) );
  CLKBUFX6 U143 ( .A(TEMP_H[48]), .Y(n110) );
  CLKINVX2 U144 ( .A(n108), .Y(n102) );
  CLKBUFX6 U145 ( .A(TEMP_H[40]), .Y(n108) );
  CLKINVX3 U146 ( .A(n121), .Y(n103) );
  INVX6 U147 ( .A(n179), .Y(n121) );
  CLKINVX4 U148 ( .A(n118), .Y(n111) );
  INVX6 U149 ( .A(n215), .Y(n118) );
  CLKINVX4 U150 ( .A(n120), .Y(n112) );
  INVX6 U151 ( .A(n197), .Y(n120) );
  CLKINVX4 U152 ( .A(n117), .Y(n113) );
  INVX6 U153 ( .A(n191), .Y(n117) );
  CLKINVX4 U154 ( .A(n122), .Y(n114) );
  INVX6 U155 ( .A(n209), .Y(n122) );
  CLKINVX4 U156 ( .A(n119), .Y(n115) );
  INVX6 U157 ( .A(n185), .Y(n119) );
  CLKINVX4 U158 ( .A(n123), .Y(n116) );
  INVX6 U159 ( .A(n203), .Y(n123) );
  OAI22X1 U160 ( .A0(n75), .A1(n655), .B0(n654), .B1(n653), .Y(
        MULi_1_mult_15_n78) );
  NAND2X2 U161 ( .A(n151), .B(n188), .Y(n183) );
  NAND2X2 U162 ( .A(n152), .B(n218), .Y(n213) );
  NAND2X2 U163 ( .A(n154), .B(n194), .Y(n189) );
  NAND2X2 U164 ( .A(n148), .B(n212), .Y(n207) );
  NAND2X2 U165 ( .A(n153), .B(n200), .Y(n195) );
  NAND2X2 U166 ( .A(n149), .B(n206), .Y(n201) );
  NAND2X2 U167 ( .A(n150), .B(n182), .Y(n177) );
  AOI22X2 U168 ( .A0(n420), .A1(n404), .B0(n85), .B1(n151), .Y(n405) );
  AOI22X2 U169 ( .A0(n420), .A1(n402), .B0(n91), .B1(n151), .Y(n403) );
  AOI22X2 U170 ( .A0(n676), .A1(n658), .B0(n92), .B1(n148), .Y(n659) );
  AOI22X2 U171 ( .A0(n676), .A1(n660), .B0(n84), .B1(n148), .Y(n661) );
  AOI22X2 U172 ( .A0(n484), .A1(n464), .B0(TEMP_H[23]), .B1(n154), .Y(n465) );
  NOR2X2 U173 ( .A(n149), .B(n235), .Y(n226) );
  AOI22X2 U174 ( .A0(n612), .A1(n596), .B0(n82), .B1(n153), .Y(n597) );
  AOI22X2 U175 ( .A0(n292), .A1(n272), .B0(TEMP_H[55]), .B1(n149), .Y(n273) );
  NOR2X2 U176 ( .A(n153), .B(n555), .Y(n224) );
  AOI22X2 U177 ( .A0(n292), .A1(n276), .B0(n86), .B1(n149), .Y(n277) );
  AOI22X2 U178 ( .A0(n612), .A1(n594), .B0(n90), .B1(n153), .Y(n595) );
  AOI22X2 U179 ( .A0(n612), .A1(n592), .B0(TEMP_H[39]), .B1(n153), .Y(n593) );
  AOI22X2 U180 ( .A0(n484), .A1(n466), .B0(n89), .B1(n154), .Y(n467) );
  AOI22X2 U181 ( .A0(n292), .A1(n274), .B0(n94), .B1(n149), .Y(n275) );
  NOR2X2 U182 ( .A(n154), .B(n427), .Y(n222) );
  AOI22X2 U183 ( .A0(n484), .A1(n468), .B0(n83), .B1(n154), .Y(n469) );
  AOI22X2 U184 ( .A0(n548), .A1(n532), .B0(n81), .B1(n152), .Y(n533) );
  NOR2X2 U185 ( .A(n150), .B(n299), .Y(n232) );
  NOR2X2 U186 ( .A(n151), .B(n363), .Y(n220) );
  AOI22X2 U187 ( .A0(n548), .A1(n530), .B0(n88), .B1(n152), .Y(n531) );
  NOR2X2 U188 ( .A(n152), .B(n491), .Y(n230) );
  AOI22X2 U189 ( .A0(n356), .A1(n340), .B0(n87), .B1(n150), .Y(n341) );
  AOI22X2 U190 ( .A0(n676), .A1(n656), .B0(TEMP_H[47]), .B1(n148), .Y(n657) );
  AOI22X2 U191 ( .A0(n356), .A1(n336), .B0(TEMP_H[7]), .B1(n150), .Y(n337) );
  AOI22X2 U192 ( .A0(n356), .A1(n342), .B0(TEMP_H[4]), .B1(n150), .Y(n343) );
  NOR2X2 U193 ( .A(n148), .B(n619), .Y(n228) );
  AOI22X2 U194 ( .A0(n548), .A1(n528), .B0(TEMP_H[31]), .B1(n152), .Y(n529) );
  AOI22X2 U195 ( .A0(n420), .A1(n400), .B0(TEMP_H[15]), .B1(n151), .Y(n401) );
  INVX16 U196 ( .A(n612), .Y(n153) );
  INVX16 U197 ( .A(n420), .Y(n151) );
  INVX16 U198 ( .A(n548), .Y(n152) );
  INVX16 U199 ( .A(n292), .Y(n149) );
  INVX16 U200 ( .A(n356), .Y(n150) );
  INVX16 U201 ( .A(n484), .Y(n154) );
  INVX16 U202 ( .A(n676), .Y(n148) );
  BUFX12 U203 ( .A(SR_to_MUL[33]), .Y(n612) );
  BUFX12 U204 ( .A(SR_to_MUL[49]), .Y(n292) );
  BUFX10 U205 ( .A(SR_to_MUL[55]), .Y(n289) );
  BUFX10 U206 ( .A(SR_to_MUL[31]), .Y(n545) );
  BUFX10 U207 ( .A(SR_to_MUL[39]), .Y(n609) );
  BUFX10 U208 ( .A(SR_to_MUL[47]), .Y(n673) );
  BUFX12 U209 ( .A(SR_to_MUL[9]), .Y(n420) );
  BUFX12 U210 ( .A(SR_to_MUL[7]), .Y(n353) );
  BUFX12 U211 ( .A(SR_to_MUL[25]), .Y(n548) );
  BUFX10 U212 ( .A(SR_to_MUL[1]), .Y(n356) );
  BUFX10 U213 ( .A(SR_to_MUL[23]), .Y(n481) );
  BUFX12 U214 ( .A(SR_to_MUL[17]), .Y(n484) );
  BUFX12 U215 ( .A(SR_to_MUL[41]), .Y(n676) );
  BUFX10 U216 ( .A(SR_to_MUL[15]), .Y(n417) );
  INVX2 U217 ( .A(MULi_5_mult_15_n1), .Y(MUL_to_PIPE1[31]) );
  INVX2 U218 ( .A(MULi_1_mult_15_n1), .Y(MUL_to_PIPE1[95]) );
  INVX2 U219 ( .A(MULi_0_mult_15_n1), .Y(MUL_to_PIPE1[111]) );
  INVX2 U220 ( .A(MULi_4_mult_15_n1), .Y(MUL_to_PIPE1[47]) );
  INVX2 U221 ( .A(MULi_3_mult_15_n1), .Y(MUL_to_PIPE1[63]) );
  INVX2 U222 ( .A(MULi_2_mult_15_n1), .Y(MUL_to_PIPE1[79]) );
  INVX2 U223 ( .A(MULi_6_mult_15_n1), .Y(MUL_to_PIPE1[15]) );
  INVX2 U224 ( .A(ADD2_1_add_16_DP_OP_277_5600_1_n1), .Y(ADD_esteso_10__17_)
         );
  INVX2 U225 ( .A(ADD2_2_add_16_DP_OP_276_702_2_n1), .Y(ADD_esteso_11__17_) );
  OAI22X1 U226 ( .A0(n75), .A1(n650), .B0(n654), .B1(n651), .Y(
        MULi_1_mult_15_n76) );
  OAI22X1 U227 ( .A0(n78), .A1(n458), .B0(n462), .B1(n459), .Y(
        MULi_4_mult_15_n76) );
  OAI22X1 U228 ( .A0(n75), .A1(n651), .B0(n654), .B1(n655), .Y(
        MULi_1_mult_15_n77) );
  INVX2 U229 ( .A(n168), .Y(n169) );
  INVX2 U230 ( .A(n158), .Y(n159) );
  OAI2BB2X2 U231 ( .B0(n690), .B1(n689), .A0N(ADD_esteso_13__9_), .A1N(
        ADD_esteso_12__9_), .Y(ADD3_1_add_16_carry_10_) );
  OAI22X1 U232 ( .A0(n77), .A1(n586), .B0(n590), .B1(n587), .Y(
        MULi_2_mult_15_n76) );
  INVX2 U233 ( .A(n166), .Y(n167) );
  INVX2 U234 ( .A(n160), .Y(n161) );
  OAI22X1 U235 ( .A0(n79), .A1(n395), .B0(n398), .B1(n399), .Y(
        MULi_5_mult_15_n77) );
  INVX2 U236 ( .A(n164), .Y(n165) );
  INVX2 U237 ( .A(n162), .Y(n163) );
  AOI222X2 U238 ( .A0(ADD_esteso_12__8_), .A1(ADD_esteso_13__8_), .B0(
        ADD_esteso_12__8_), .B1(n688), .C0(ADD_esteso_13__8_), .C1(n688), .Y(
        n690) );
  AO22X2 U239 ( .A0(n455), .A1(n453), .B0(n428), .B1(n170), .Y(n158) );
  AO22X2 U240 ( .A0(n583), .A1(n581), .B0(n556), .B1(n173), .Y(n164) );
  AO22X2 U241 ( .A0(n519), .A1(n517), .B0(n492), .B1(n171), .Y(n160) );
  AO22X2 U242 ( .A0(n263), .A1(n261), .B0(n236), .B1(n174), .Y(n166) );
  AO22X2 U243 ( .A0(n391), .A1(n389), .B0(n364), .B1(n172), .Y(n162) );
  INVX2 U244 ( .A(n156), .Y(n157) );
  AO22X2 U245 ( .A0(n647), .A1(n645), .B0(n620), .B1(n175), .Y(n168) );
  AO22X2 U246 ( .A0(n327), .A1(n325), .B0(n300), .B1(n176), .Y(n156) );
  BUFX3 U247 ( .A(n390), .Y(n172) );
  BUFX3 U248 ( .A(n518), .Y(n171) );
  BUFX3 U249 ( .A(n582), .Y(n173) );
  BUFX3 U250 ( .A(n262), .Y(n174) );
  BUFX3 U251 ( .A(n646), .Y(n175) );
  BUFX3 U252 ( .A(n454), .Y(n170) );
  NAND2X2 U253 ( .A(n207), .B(n208), .Y(n621) );
  NAND2X2 U254 ( .A(n177), .B(n178), .Y(n301) );
  NAND2X2 U255 ( .A(n183), .B(n184), .Y(n365) );
  NAND2X2 U256 ( .A(n213), .B(n214), .Y(n493) );
  NAND2X2 U257 ( .A(n195), .B(n196), .Y(n557) );
  NAND2X2 U258 ( .A(n201), .B(n202), .Y(n237) );
  NAND2X2 U259 ( .A(n189), .B(n190), .Y(n429) );
  NOR2X2 U260 ( .A(n78), .B(n479), .Y(MULi_4_mult_15_n79) );
  NOR2X2 U261 ( .A(n76), .B(n287), .Y(MULi_0_mult_15_n79) );
  NOR2X2 U262 ( .A(n74), .B(n543), .Y(MULi_3_mult_15_n79) );
  NOR2X2 U263 ( .A(n75), .B(n671), .Y(MULi_1_mult_15_n79) );
  NOR2X2 U264 ( .A(n79), .B(n415), .Y(MULi_5_mult_15_n79) );
  INVX2 U265 ( .A(MULi_1_mult_15_n21), .Y(MULi_1_mult_15_n22) );
  INVX2 U266 ( .A(MULi_5_mult_15_n21), .Y(MULi_5_mult_15_n22) );
  NOR2X2 U267 ( .A(n77), .B(n607), .Y(MULi_2_mult_15_n79) );
  INVX2 U268 ( .A(MULi_5_mult_15_n15), .Y(MULi_5_mult_15_n16) );
  INVX2 U269 ( .A(MULi_1_mult_15_n15), .Y(MULi_1_mult_15_n16) );
  INVX2 U270 ( .A(MULi_4_mult_15_n21), .Y(MULi_4_mult_15_n22) );
  ADDHX1 U271 ( .A(MULi_3_mult_15_n81), .B(MULi_3_mult_15_n52), .CO(
        MULi_3_mult_15_n39), .S(MULi_3_mult_15_n40) );
  INVX2 U272 ( .A(MULi_0_mult_15_n15), .Y(MULi_0_mult_15_n16) );
  INVX2 U273 ( .A(MULi_4_mult_15_n15), .Y(MULi_4_mult_15_n16) );
  NOR2X2 U274 ( .A(n80), .B(n351), .Y(MULi_6_mult_15_n79) );
  ADDHX1 U275 ( .A(MULi_6_mult_15_n81), .B(MULi_6_mult_15_n52), .CO(
        MULi_6_mult_15_n39), .S(MULi_6_mult_15_n40) );
  INVX2 U276 ( .A(MULi_0_mult_15_n21), .Y(MULi_0_mult_15_n22) );
  ADDHX1 U277 ( .A(MULi_0_mult_15_n81), .B(MULi_0_mult_15_n52), .CO(
        MULi_0_mult_15_n39), .S(MULi_0_mult_15_n40) );
  INVX4 U278 ( .A(n80), .Y(n327) );
  INVX2 U279 ( .A(MULi_2_mult_15_n21), .Y(MULi_2_mult_15_n22) );
  ADDHX1 U280 ( .A(MULi_2_mult_15_n81), .B(MULi_2_mult_15_n52), .CO(
        MULi_2_mult_15_n39), .S(MULi_2_mult_15_n40) );
  ADDHX1 U281 ( .A(MULi_1_mult_15_n81), .B(MULi_1_mult_15_n52), .CO(
        MULi_1_mult_15_n39), .S(MULi_1_mult_15_n40) );
  INVX2 U282 ( .A(MULi_2_mult_15_n15), .Y(MULi_2_mult_15_n16) );
  INVX2 U283 ( .A(MULi_3_mult_15_n21), .Y(MULi_3_mult_15_n22) );
  ADDHX1 U284 ( .A(MULi_5_mult_15_n81), .B(MULi_5_mult_15_n52), .CO(
        MULi_5_mult_15_n39), .S(MULi_5_mult_15_n40) );
  INVX2 U285 ( .A(MULi_6_mult_15_n15), .Y(MULi_6_mult_15_n16) );
  INVX2 U286 ( .A(MULi_6_mult_15_n21), .Y(MULi_6_mult_15_n22) );
  INVX2 U287 ( .A(MULi_3_mult_15_n15), .Y(MULi_3_mult_15_n16) );
  ADDHX1 U288 ( .A(MULi_4_mult_15_n81), .B(MULi_4_mult_15_n52), .CO(
        MULi_4_mult_15_n39), .S(MULi_4_mult_15_n40) );
  AO21X2 U289 ( .A0(n615), .A1(n616), .B0(n570), .Y(MULi_2_mult_15_n64) );
  NOR2X2 U290 ( .A(n415), .B(n421), .Y(MULi_5_mult_15_n63) );
  AOI222X2 U291 ( .A0(ADD_esteso_12__4_), .A1(ADD_esteso_13__4_), .B0(
        ADD_esteso_12__4_), .B1(n684), .C0(ADD_esteso_13__4_), .C1(n684), .Y(
        n685) );
  NOR2X2 U292 ( .A(n543), .B(n549), .Y(MULi_3_mult_15_n63) );
  AO21X2 U293 ( .A0(n613), .A1(n614), .B0(n559), .Y(MULi_2_mult_15_n56) );
  NOR2X2 U294 ( .A(n423), .B(n415), .Y(MULi_5_mult_15_n71) );
  AO21X2 U295 ( .A0(n421), .A1(n422), .B0(n367), .Y(MULi_5_mult_15_n56) );
  AO21X2 U296 ( .A0(n423), .A1(n424), .B0(n378), .Y(MULi_5_mult_15_n64) );
  NOR2X2 U297 ( .A(n551), .B(n543), .Y(MULi_3_mult_15_n71) );
  NOR2X2 U298 ( .A(n607), .B(n613), .Y(MULi_2_mult_15_n63) );
  AO21X2 U299 ( .A0(n293), .A1(n294), .B0(n239), .Y(MULi_0_mult_15_n56) );
  AO21X2 U300 ( .A0(n295), .A1(n296), .B0(n250), .Y(MULi_0_mult_15_n64) );
  NOR2X2 U301 ( .A(n359), .B(n351), .Y(MULi_6_mult_15_n71) );
  NOR2X2 U302 ( .A(n351), .B(n357), .Y(MULi_6_mult_15_n63) );
  AO21X2 U303 ( .A0(n485), .A1(n486), .B0(n431), .Y(MULi_4_mult_15_n56) );
  AO21X2 U304 ( .A0(n487), .A1(n488), .B0(n442), .Y(MULi_4_mult_15_n64) );
  NOR2X2 U305 ( .A(n671), .B(n677), .Y(MULi_1_mult_15_n63) );
  AO21X2 U306 ( .A0(n679), .A1(n680), .B0(n634), .Y(MULi_1_mult_15_n64) );
  NOR2X2 U307 ( .A(n679), .B(n671), .Y(MULi_1_mult_15_n71) );
  AO21X2 U308 ( .A0(n677), .A1(n678), .B0(n623), .Y(MULi_1_mult_15_n56) );
  NOR2X2 U309 ( .A(n479), .B(n485), .Y(MULi_4_mult_15_n63) );
  NOR2X2 U310 ( .A(n487), .B(n479), .Y(MULi_4_mult_15_n71) );
  AO21X2 U311 ( .A0(n359), .A1(n360), .B0(n314), .Y(MULi_6_mult_15_n64) );
  AO21X2 U312 ( .A0(n357), .A1(n358), .B0(n303), .Y(MULi_6_mult_15_n56) );
  NOR2X2 U313 ( .A(n295), .B(n287), .Y(MULi_0_mult_15_n71) );
  NOR2X2 U314 ( .A(n615), .B(n607), .Y(MULi_2_mult_15_n71) );
  AO21X2 U315 ( .A0(n551), .A1(n552), .B0(n506), .Y(MULi_3_mult_15_n64) );
  AO21X2 U316 ( .A0(n549), .A1(n550), .B0(n495), .Y(MULi_3_mult_15_n56) );
  NOR2X2 U317 ( .A(n287), .B(n293), .Y(MULi_0_mult_15_n63) );
  BUFX8 U318 ( .A(n516), .Y(n551) );
  NAND2X2 U319 ( .A(n292), .B(n205), .Y(n202) );
  AND2X2 U320 ( .A(n203), .B(n204), .Y(n206) );
  BUFX8 U321 ( .A(n324), .Y(n359) );
  BUFX8 U322 ( .A(n322), .Y(n360) );
  NAND2X2 U323 ( .A(n676), .B(n211), .Y(n208) );
  BUFX8 U324 ( .A(n452), .Y(n487) );
  BUFX8 U325 ( .A(n450), .Y(n488) );
  BUFX8 U326 ( .A(n313), .Y(n357) );
  BUFX8 U327 ( .A(n375), .Y(n422) );
  BUFX8 U328 ( .A(n441), .Y(n485) );
  AND2X2 U329 ( .A(n185), .B(n186), .Y(n188) );
  BUFX8 U330 ( .A(n439), .Y(n486) );
  AND2X2 U331 ( .A(n209), .B(n210), .Y(n212) );
  NAND2X2 U332 ( .A(n420), .B(n187), .Y(n184) );
  BUFX8 U333 ( .A(n311), .Y(n358) );
  BUFX8 U334 ( .A(n247), .Y(n294) );
  AND2X2 U335 ( .A(n197), .B(n198), .Y(n200) );
  BUFX8 U336 ( .A(n249), .Y(n293) );
  BUFX8 U337 ( .A(n386), .Y(n424) );
  BUFX8 U338 ( .A(n580), .Y(n615) );
  BUFX8 U339 ( .A(n258), .Y(n296) );
  BUFX8 U340 ( .A(n578), .Y(n616) );
  NAND2X2 U341 ( .A(n612), .B(n199), .Y(n196) );
  BUFX8 U342 ( .A(n631), .Y(n678) );
  BUFX8 U343 ( .A(n260), .Y(n295) );
  BUFX8 U344 ( .A(n388), .Y(n423) );
  BUFX8 U345 ( .A(n633), .Y(n677) );
  BUFX8 U346 ( .A(n503), .Y(n550) );
  NAND2X2 U347 ( .A(n356), .B(n181), .Y(n178) );
  AND2X2 U348 ( .A(n179), .B(n180), .Y(n182) );
  AND2X2 U349 ( .A(n215), .B(n216), .Y(n218) );
  BUFX8 U350 ( .A(n505), .Y(n549) );
  AND2X2 U351 ( .A(n191), .B(n192), .Y(n194) );
  NAND2X2 U352 ( .A(n548), .B(n217), .Y(n214) );
  NAND2X2 U353 ( .A(n484), .B(n193), .Y(n190) );
  BUFX8 U354 ( .A(n567), .Y(n614) );
  BUFX8 U355 ( .A(n569), .Y(n613) );
  BUFX8 U356 ( .A(n644), .Y(n679) );
  BUFX8 U357 ( .A(n514), .Y(n552) );
  BUFX8 U358 ( .A(n642), .Y(n680) );
  BUFX8 U359 ( .A(n377), .Y(n421) );
  AOI22X2 U360 ( .A0(n675), .A1(n618), .B0(SR_to_MUL[44]), .B1(n652), .Y(n644)
         );
  AOI33X2 U361 ( .A0(n419), .A1(SR_to_MUL[12]), .A2(n384), .B0(n418), .B1(n362), .B2(n396), .Y(n386) );
  AOI33X2 U362 ( .A0(n675), .A1(SR_to_MUL[44]), .A2(n640), .B0(n674), .B1(n618), .B2(n652), .Y(n642) );
  AOI22X2 U363 ( .A0(n675), .A1(n671), .B0(TEMP_H[40]), .B1(n652), .Y(n653) );
  INVX2 U364 ( .A(n480), .Y(n191) );
  AOI22X2 U365 ( .A0(n674), .A1(n671), .B0(TEMP_H[40]), .B1(n640), .Y(n641) );
  INVX2 U366 ( .A(n352), .Y(n179) );
  AOI22X2 U367 ( .A0(n105), .A1(n437), .B0(n481), .B1(n96), .Y(n438) );
  AOI33X2 U368 ( .A0(n290), .A1(SR_to_MUL[54]), .A2(n245), .B0(n289), .B1(n233), .B2(n256), .Y(n247) );
  AOI22X2 U369 ( .A0(n418), .A1(n415), .B0(TEMP_H[8]), .B1(n384), .Y(n385) );
  AOI22X2 U370 ( .A0(n674), .A1(n617), .B0(SR_to_MUL[46]), .B1(n640), .Y(n633)
         );
  AOI22X2 U371 ( .A0(n290), .A1(n233), .B0(SR_to_MUL[54]), .B1(n256), .Y(n249)
         );
  AOI22X2 U372 ( .A0(n291), .A1(n234), .B0(SR_to_MUL[52]), .B1(n268), .Y(n260)
         );
  AOI22X2 U373 ( .A0(n419), .A1(n362), .B0(SR_to_MUL[12]), .B1(n396), .Y(n388)
         );
  AOI33X2 U374 ( .A0(n674), .A1(SR_to_MUL[46]), .A2(n629), .B0(n673), .B1(n617), .B2(n640), .Y(n631) );
  AOI33X2 U375 ( .A0(n291), .A1(SR_to_MUL[52]), .A2(n256), .B0(n290), .B1(n234), .B2(n268), .Y(n258) );
  AOI22X2 U376 ( .A0(n482), .A1(n479), .B0(TEMP_H[16]), .B1(n448), .Y(n449) );
  AOI22X2 U377 ( .A0(n483), .A1(n479), .B0(TEMP_H[16]), .B1(n460), .Y(n461) );
  AOI22X2 U378 ( .A0(n419), .A1(n415), .B0(TEMP_H[8]), .B1(n396), .Y(n397) );
  AOI22X2 U379 ( .A0(n355), .A1(n351), .B0(TEMP_H[0]), .B1(n332), .Y(n333) );
  AOI22X2 U380 ( .A0(n354), .A1(n351), .B0(TEMP_H[0]), .B1(n320), .Y(n321) );
  AOI33X2 U381 ( .A0(n354), .A1(SR_to_MUL[6]), .A2(n309), .B0(n353), .B1(n297), 
        .B2(n320), .Y(n311) );
  AOI22X2 U382 ( .A0(n291), .A1(n287), .B0(TEMP_H[48]), .B1(n268), .Y(n269) );
  INVX2 U383 ( .A(n672), .Y(n209) );
  AOI33X2 U384 ( .A0(n418), .A1(SR_to_MUL[14]), .A2(n373), .B0(n417), .B1(n361), .B2(n384), .Y(n375) );
  AOI33X2 U385 ( .A0(n482), .A1(SR_to_MUL[22]), .A2(n437), .B0(n481), .B1(n425), .B2(n448), .Y(n439) );
  AOI22X2 U386 ( .A0(n290), .A1(n287), .B0(TEMP_H[48]), .B1(n256), .Y(n257) );
  INVX2 U387 ( .A(n416), .Y(n185) );
  AOI22X2 U388 ( .A0(n354), .A1(n297), .B0(SR_to_MUL[6]), .B1(n320), .Y(n313)
         );
  AOI22X2 U389 ( .A0(n482), .A1(n425), .B0(SR_to_MUL[22]), .B1(n448), .Y(n441)
         );
  AOI33X2 U390 ( .A0(n483), .A1(SR_to_MUL[20]), .A2(n448), .B0(n482), .B1(n426), .B2(n460), .Y(n450) );
  NOR2X2 U391 ( .A(n120), .B(n100), .Y(MUL_to_PIPE1[64]) );
  AOI22X2 U392 ( .A0(n483), .A1(n426), .B0(SR_to_MUL[20]), .B1(n460), .Y(n452)
         );
  NOR2X2 U393 ( .A(n119), .B(n97), .Y(MUL_to_PIPE1[16]) );
  AOI22X2 U394 ( .A0(n108), .A1(n629), .B0(n673), .B1(n102), .Y(n630) );
  AOI22X2 U395 ( .A0(n110), .A1(n245), .B0(n289), .B1(n101), .Y(n246) );
  NOR2X2 U396 ( .A(n118), .B(n98), .Y(MUL_to_PIPE1[48]) );
  AOI33X2 U397 ( .A0(n355), .A1(SR_to_MUL[4]), .A2(n320), .B0(n354), .B1(n298), 
        .B2(n332), .Y(n322) );
  NOR2X2 U398 ( .A(n123), .B(n101), .Y(MUL_to_PIPE1[96]) );
  AOI22X2 U399 ( .A0(n355), .A1(n298), .B0(SR_to_MUL[4]), .B1(n332), .Y(n324)
         );
  NOR2X2 U400 ( .A(n117), .B(n96), .Y(MUL_to_PIPE1[32]) );
  AOI22X2 U401 ( .A0(n107), .A1(n373), .B0(n417), .B1(n97), .Y(n374) );
  NOR2X2 U402 ( .A(n121), .B(n99), .Y(MUL_to_PIPE1[0]) );
  AOI22X2 U403 ( .A0(n109), .A1(n309), .B0(n353), .B1(n99), .Y(n310) );
  INVX2 U404 ( .A(n288), .Y(n203) );
  NOR2X2 U405 ( .A(n122), .B(n102), .Y(MUL_to_PIPE1[80]) );
  AOI22X2 U406 ( .A0(n95), .A1(n309), .B0(n353), .B1(n342), .Y(n155) );
  AOI22X2 U407 ( .A0(n418), .A1(n361), .B0(SR_to_MUL[14]), .B1(n384), .Y(n377)
         );
  AOI33X2 U408 ( .A0(n547), .A1(SR_to_MUL[28]), .A2(n512), .B0(n546), .B1(n490), .B2(n524), .Y(n514) );
  INVX2 U409 ( .A(n608), .Y(n197) );
  AOI22X2 U410 ( .A0(n611), .A1(n607), .B0(TEMP_H[32]), .B1(n588), .Y(n589) );
  AOI22X2 U411 ( .A0(n546), .A1(n489), .B0(SR_to_MUL[30]), .B1(n512), .Y(n505)
         );
  AOI22X2 U412 ( .A0(n611), .A1(n554), .B0(SR_to_MUL[36]), .B1(n588), .Y(n580)
         );
  AOI33X2 U413 ( .A0(n611), .A1(SR_to_MUL[36]), .A2(n576), .B0(n610), .B1(n554), .B2(n588), .Y(n578) );
  AOI22X2 U414 ( .A0(n610), .A1(n607), .B0(TEMP_H[32]), .B1(n576), .Y(n577) );
  AOI22X2 U415 ( .A0(n610), .A1(n553), .B0(SR_to_MUL[38]), .B1(n576), .Y(n569)
         );
  AOI22X2 U416 ( .A0(n547), .A1(n543), .B0(TEMP_H[24]), .B1(n524), .Y(n525) );
  AOI22X2 U417 ( .A0(n106), .A1(n565), .B0(n609), .B1(n100), .Y(n566) );
  INVX2 U418 ( .A(n544), .Y(n215) );
  AOI22X2 U419 ( .A0(n547), .A1(n490), .B0(SR_to_MUL[28]), .B1(n524), .Y(n516)
         );
  AOI33X2 U420 ( .A0(n610), .A1(SR_to_MUL[38]), .A2(n565), .B0(n609), .B1(n553), .B2(n576), .Y(n567) );
  AOI33X2 U421 ( .A0(n546), .A1(SR_to_MUL[30]), .A2(n501), .B0(n545), .B1(n489), .B2(n512), .Y(n503) );
  AOI22X2 U422 ( .A0(n104), .A1(n501), .B0(n545), .B1(n98), .Y(n502) );
  AOI22X2 U423 ( .A0(n546), .A1(n543), .B0(TEMP_H[24]), .B1(n512), .Y(n513) );
  INVX12 U424 ( .A(n674), .Y(n640) );
  INVX12 U425 ( .A(n547), .Y(n524) );
  INVX12 U426 ( .A(n291), .Y(n268) );
  INVX10 U427 ( .A(n673), .Y(n629) );
  INVX10 U428 ( .A(n353), .Y(n309) );
  INVX12 U429 ( .A(n290), .Y(n256) );
  NOR2X2 U430 ( .A(SR_to_MUL[10]), .B(n420), .Y(n219) );
  NOR2X2 U431 ( .A(SR_to_MUL[2]), .B(n356), .Y(n231) );
  INVX10 U432 ( .A(n289), .Y(n245) );
  INVX10 U433 ( .A(n609), .Y(n565) );
  INVX10 U434 ( .A(n417), .Y(n373) );
  INVX12 U435 ( .A(n610), .Y(n576) );
  INVX12 U436 ( .A(n418), .Y(n384) );
  INVX12 U437 ( .A(n675), .Y(n652) );
  INVX10 U438 ( .A(n481), .Y(n437) );
  INVX12 U439 ( .A(n419), .Y(n396) );
  NOR2X2 U440 ( .A(SR_to_MUL[34]), .B(n612), .Y(n223) );
  NOR2X2 U441 ( .A(SR_to_MUL[42]), .B(n676), .Y(n227) );
  INVX12 U442 ( .A(n482), .Y(n448) );
  NOR2X2 U443 ( .A(SR_to_MUL[50]), .B(n292), .Y(n225) );
  INVX12 U444 ( .A(n611), .Y(n588) );
  INVX10 U445 ( .A(n545), .Y(n501) );
  NOR2X2 U446 ( .A(SR_to_MUL[26]), .B(n548), .Y(n229) );
  INVX12 U447 ( .A(n546), .Y(n512) );
  INVX12 U448 ( .A(n483), .Y(n460) );
  NOR2X2 U449 ( .A(SR_to_MUL[18]), .B(n484), .Y(n221) );
  INVX2 U450 ( .A(ADD_esteso_2__17_), .Y(ADD2_1_add_16_DP_OP_277_5600_1_n69)
         );
  NOR2X2 U451 ( .A(ADD_esteso_13__9_), .B(ADD_esteso_12__9_), .Y(n689) );
  OAI211X2 U452 ( .A0(ADD_esteso_13__1_), .A1(ADD_esteso_12__1_), .B0(
        ADD_esteso_12__0_), .C0(ADD_esteso_13__0_), .Y(n681) );
  INVX2 U453 ( .A(ADD_esteso_5__17_), .Y(ADD2_2_add_16_DP_OP_276_702_2_n50) );
  INVX2 U454 ( .A(ADD_esteso_6__17_), .Y(ADD2_2_add_16_DP_OP_276_702_2_n48) );
  INVX2 U455 ( .A(ADD_esteso_4__17_), .Y(ADD2_2_add_16_DP_OP_276_702_2_n49) );
  INVX2 U456 ( .A(ADD_esteso_3__17_), .Y(ADD2_1_add_16_DP_OP_277_5600_1_n66)
         );
  INVX2 U457 ( .A(ADD_esteso_1__17_), .Y(ADD2_1_add_16_DP_OP_277_5600_1_n67)
         );
  INVX2 U458 ( .A(ADD_esteso_0__17_), .Y(ADD2_1_add_16_DP_OP_277_5600_1_n68)
         );
  BUFX12 U459 ( .A(SR_to_MUL[3]), .Y(n355) );
  AOI22X4 U460 ( .A0(TEMP_H[31]), .A1(n501), .B0(n545), .B1(n528), .Y(n495) );
  AOI22X4 U461 ( .A0(TEMP_H[23]), .A1(n437), .B0(n481), .B1(n464), .Y(n431) );
  AOI22X4 U462 ( .A0(TEMP_H[39]), .A1(n565), .B0(n609), .B1(n592), .Y(n559) );
  AOI22X4 U463 ( .A0(TEMP_H[15]), .A1(n373), .B0(n417), .B1(n400), .Y(n367) );
  AOI22X4 U464 ( .A0(TEMP_H[47]), .A1(n629), .B0(n673), .B1(n656), .Y(n623) );
  AOI22X4 U465 ( .A0(TEMP_H[55]), .A1(n245), .B0(n289), .B1(n272), .Y(n239) );
  AOI22X4 U466 ( .A0(TEMP_H[31]), .A1(n512), .B0(n546), .B1(n528), .Y(n506) );
  AOI22X4 U467 ( .A0(TEMP_H[23]), .A1(n448), .B0(n482), .B1(n464), .Y(n442) );
  AOI22X4 U468 ( .A0(TEMP_H[39]), .A1(n576), .B0(n610), .B1(n592), .Y(n570) );
  AOI22X4 U469 ( .A0(TEMP_H[15]), .A1(n384), .B0(n418), .B1(n400), .Y(n378) );
  AOI22X4 U470 ( .A0(TEMP_H[47]), .A1(n640), .B0(n674), .B1(n656), .Y(n634) );
  AOI22X4 U471 ( .A0(TEMP_H[55]), .A1(n256), .B0(n290), .B1(n272), .Y(n250) );
  AOI22X4 U472 ( .A0(TEMP_H[22]), .A1(n437), .B0(n481), .B1(n466), .Y(n432) );
  AOI22X4 U473 ( .A0(TEMP_H[30]), .A1(n501), .B0(n545), .B1(n530), .Y(n496) );
  AOI22X4 U474 ( .A0(TEMP_H[14]), .A1(n373), .B0(n417), .B1(n402), .Y(n368) );
  AOI22X4 U475 ( .A0(TEMP_H[38]), .A1(n565), .B0(n609), .B1(n594), .Y(n560) );
  AOI22X4 U476 ( .A0(TEMP_H[54]), .A1(n245), .B0(n289), .B1(n274), .Y(n240) );
  AOI22X4 U477 ( .A0(TEMP_H[46]), .A1(n629), .B0(n673), .B1(n658), .Y(n624) );
  OAI32X4 U478 ( .A0(n437), .A1(n105), .A2(n485), .B0(n486), .B1(n437), .Y(
        MULi_4_mult_15_n52) );
  OAI32X4 U479 ( .A0(n501), .A1(n104), .A2(n549), .B0(n550), .B1(n501), .Y(
        MULi_3_mult_15_n52) );
  OAI32X4 U480 ( .A0(n373), .A1(n107), .A2(n421), .B0(n422), .B1(n373), .Y(
        MULi_5_mult_15_n52) );
  OAI32X4 U481 ( .A0(n565), .A1(n106), .A2(n613), .B0(n614), .B1(n565), .Y(
        MULi_2_mult_15_n52) );
  OAI32X4 U482 ( .A0(n309), .A1(n109), .A2(n357), .B0(n358), .B1(n309), .Y(
        MULi_6_mult_15_n52) );
  OAI32X4 U483 ( .A0(n629), .A1(n108), .A2(n677), .B0(n678), .B1(n629), .Y(
        MULi_1_mult_15_n52) );
  OAI32X4 U484 ( .A0(n245), .A1(n110), .A2(n293), .B0(n294), .B1(n245), .Y(
        MULi_0_mult_15_n52) );
  AOI22X4 U485 ( .A0(TEMP_H[7]), .A1(n309), .B0(n353), .B1(n336), .Y(n303) );
  AOI22X4 U486 ( .A0(n483), .A1(n475), .B0(TEMP_H[17]), .B1(n460), .Y(n463) );
  AOI22X4 U487 ( .A0(n547), .A1(n539), .B0(TEMP_H[25]), .B1(n524), .Y(n527) );
  AOI22X4 U488 ( .A0(n419), .A1(n411), .B0(TEMP_H[9]), .B1(n396), .Y(n399) );
  AOI22X4 U489 ( .A0(n611), .A1(n603), .B0(TEMP_H[33]), .B1(n588), .Y(n591) );
  AOI22X4 U490 ( .A0(n355), .A1(n347), .B0(TEMP_H[1]), .B1(n332), .Y(n335) );
  INVX12 U491 ( .A(n355), .Y(n332) );
  AOI22X4 U492 ( .A0(n675), .A1(n667), .B0(TEMP_H[41]), .B1(n652), .Y(n655) );
  AOI22X4 U493 ( .A0(n291), .A1(n283), .B0(TEMP_H[49]), .B1(n268), .Y(n271) );
  AOI22X4 U494 ( .A0(TEMP_H[6]), .A1(n309), .B0(n353), .B1(n338), .Y(n304) );
  ADDHX2 U495 ( .A(MULi_6_mult_15_n83), .B(MULi_6_mult_15_n53), .CO(
        MULi_6_mult_15_n46), .S(MULi_6_mult_15_n47) );
  OAI32X4 U496 ( .A0(SR_to_MUL[0]), .A1(TEMP_H[4]), .A2(n150), .B0(n341), .B1(
        n121), .Y(MULi_6_mult_15_n83) );
  ADDHX2 U497 ( .A(MULi_3_mult_15_n83), .B(MULi_3_mult_15_n53), .CO(
        MULi_3_mult_15_n46), .S(MULi_3_mult_15_n47) );
  OAI32X4 U498 ( .A0(SR_to_MUL[24]), .A1(TEMP_H[28]), .A2(n152), .B0(n533), 
        .B1(n118), .Y(MULi_3_mult_15_n83) );
  ADDHX2 U499 ( .A(MULi_4_mult_15_n83), .B(MULi_4_mult_15_n53), .CO(
        MULi_4_mult_15_n46), .S(MULi_4_mult_15_n47) );
  OAI32X4 U500 ( .A0(SR_to_MUL[16]), .A1(TEMP_H[20]), .A2(n154), .B0(n469), 
        .B1(n117), .Y(MULi_4_mult_15_n83) );
  ADDHX2 U501 ( .A(MULi_2_mult_15_n83), .B(MULi_2_mult_15_n53), .CO(
        MULi_2_mult_15_n46), .S(MULi_2_mult_15_n47) );
  OAI32X4 U502 ( .A0(SR_to_MUL[32]), .A1(TEMP_H[36]), .A2(n153), .B0(n597), 
        .B1(n120), .Y(MULi_2_mult_15_n83) );
  ADDHX2 U503 ( .A(MULi_5_mult_15_n83), .B(MULi_5_mult_15_n53), .CO(
        MULi_5_mult_15_n46), .S(MULi_5_mult_15_n47) );
  OAI32X4 U504 ( .A0(SR_to_MUL[8]), .A1(TEMP_H[12]), .A2(n151), .B0(n405), 
        .B1(n119), .Y(MULi_5_mult_15_n83) );
  ADDHX2 U505 ( .A(MULi_1_mult_15_n83), .B(MULi_1_mult_15_n53), .CO(
        MULi_1_mult_15_n46), .S(MULi_1_mult_15_n47) );
  OAI32X4 U506 ( .A0(SR_to_MUL[40]), .A1(TEMP_H[44]), .A2(n148), .B0(n661), 
        .B1(n122), .Y(MULi_1_mult_15_n83) );
  ADDHX2 U507 ( .A(MULi_0_mult_15_n83), .B(MULi_0_mult_15_n53), .CO(
        MULi_0_mult_15_n46), .S(MULi_0_mult_15_n47) );
  OAI32X4 U508 ( .A0(SR_to_MUL[48]), .A1(TEMP_H[52]), .A2(n149), .B0(n277), 
        .B1(n123), .Y(MULi_0_mult_15_n83) );
  AOI222X2 U509 ( .A0(ADD_esteso_12__6_), .A1(ADD_esteso_13__6_), .B0(
        ADD_esteso_12__6_), .B1(n686), .C0(ADD_esteso_13__6_), .C1(n686), .Y(
        n687) );
  AOI222X2 U510 ( .A0(ADD_esteso_12__2_), .A1(ADD_esteso_13__2_), .B0(
        ADD_esteso_12__2_), .B1(n682), .C0(ADD_esteso_13__2_), .C1(n682), .Y(
        n683) );
  OAI22X4 U511 ( .A0(n359), .A1(n314), .B0(n360), .B1(n315), .Y(
        MULi_6_mult_15_n21) );
  AOI221X2 U512 ( .A0(SR_to_MUL[18]), .A1(n483), .B0(n427), .B1(n460), .C0(
        n455), .Y(n454) );
  AOI221X2 U513 ( .A0(SR_to_MUL[26]), .A1(n547), .B0(n491), .B1(n524), .C0(
        n519), .Y(n518) );
  AOI221X2 U514 ( .A0(SR_to_MUL[10]), .A1(n419), .B0(n363), .B1(n396), .C0(
        n391), .Y(n390) );
  AOI221X2 U515 ( .A0(SR_to_MUL[34]), .A1(n611), .B0(n555), .B1(n588), .C0(
        n583), .Y(n582) );
  AOI221X2 U516 ( .A0(SR_to_MUL[50]), .A1(n291), .B0(n235), .B1(n268), .C0(
        n263), .Y(n262) );
  AOI221X2 U517 ( .A0(SR_to_MUL[42]), .A1(n675), .B0(n619), .B1(n652), .C0(
        n647), .Y(n646) );
  AOI221X4 U518 ( .A0(SR_to_MUL[2]), .A1(n355), .B0(n299), .B1(n332), .C0(n327), .Y(n176) );
  AOI221X2 U519 ( .A0(SR_to_MUL[2]), .A1(n355), .B0(n299), .B1(n332), .C0(n327), .Y(n326) );
  NAND2X2 U520 ( .A(n430), .B(n429), .Y(MULi_4_mult_15_n34) );
  AOI2BB2X4 U521 ( .B0(n455), .B1(n428), .A0N(n462), .A1N(n456), .Y(n430) );
  NAND2X2 U522 ( .A(n366), .B(n365), .Y(MULi_5_mult_15_n34) );
  AOI2BB2X4 U523 ( .B0(n391), .B1(n364), .A0N(n398), .A1N(n392), .Y(n366) );
  NAND2X2 U524 ( .A(n494), .B(n493), .Y(MULi_3_mult_15_n34) );
  AOI2BB2X4 U525 ( .B0(n519), .B1(n492), .A0N(n526), .A1N(n520), .Y(n494) );
  NAND2X2 U526 ( .A(n302), .B(n301), .Y(MULi_6_mult_15_n34) );
  AOI2BB2X4 U527 ( .B0(n327), .B1(n300), .A0N(n334), .A1N(n328), .Y(n302) );
  NAND2X2 U528 ( .A(n558), .B(n557), .Y(MULi_2_mult_15_n34) );
  AOI2BB2X4 U529 ( .B0(n583), .B1(n556), .A0N(n590), .A1N(n584), .Y(n558) );
  NAND2X2 U530 ( .A(n238), .B(n237), .Y(MULi_0_mult_15_n34) );
  AOI2BB2X4 U531 ( .B0(n263), .B1(n236), .A0N(n270), .A1N(n264), .Y(n238) );
  NAND2X2 U532 ( .A(n622), .B(n621), .Y(MULi_1_mult_15_n34) );
  AOI2BB2X4 U533 ( .B0(n647), .B1(n620), .A0N(n654), .A1N(n648), .Y(n622) );
  OAI32X4 U534 ( .A0(SR_to_MUL[16]), .A1(TEMP_H[18]), .A2(n154), .B0(n473), 
        .B1(n480), .Y(MULi_4_mult_15_n85) );
  OAI32X4 U535 ( .A0(SR_to_MUL[16]), .A1(TEMP_H[19]), .A2(n154), .B0(n471), 
        .B1(n117), .Y(MULi_4_mult_15_n84) );
  OAI32X4 U536 ( .A0(SR_to_MUL[24]), .A1(TEMP_H[26]), .A2(n152), .B0(n537), 
        .B1(n544), .Y(MULi_3_mult_15_n85) );
  OAI32X4 U537 ( .A0(SR_to_MUL[24]), .A1(TEMP_H[27]), .A2(n152), .B0(n535), 
        .B1(n118), .Y(MULi_3_mult_15_n84) );
  OAI32X4 U538 ( .A0(SR_to_MUL[8]), .A1(TEMP_H[10]), .A2(n151), .B0(n409), 
        .B1(n416), .Y(MULi_5_mult_15_n85) );
  OAI32X4 U539 ( .A0(SR_to_MUL[8]), .A1(TEMP_H[11]), .A2(n151), .B0(n407), 
        .B1(n119), .Y(MULi_5_mult_15_n84) );
  OAI32X4 U540 ( .A0(SR_to_MUL[32]), .A1(TEMP_H[34]), .A2(n153), .B0(n601), 
        .B1(n608), .Y(MULi_2_mult_15_n85) );
  OAI32X4 U541 ( .A0(SR_to_MUL[32]), .A1(TEMP_H[35]), .A2(n153), .B0(n599), 
        .B1(n120), .Y(MULi_2_mult_15_n84) );
  OAI32X4 U542 ( .A0(SR_to_MUL[0]), .A1(TEMP_H[2]), .A2(n150), .B0(n345), .B1(
        n352), .Y(MULi_6_mult_15_n85) );
  OAI32X4 U543 ( .A0(SR_to_MUL[0]), .A1(TEMP_H[3]), .A2(n150), .B0(n343), .B1(
        n121), .Y(MULi_6_mult_15_n84) );
  OAI32X4 U544 ( .A0(SR_to_MUL[40]), .A1(TEMP_H[42]), .A2(n148), .B0(n665), 
        .B1(n672), .Y(MULi_1_mult_15_n85) );
  OAI32X4 U545 ( .A0(SR_to_MUL[40]), .A1(TEMP_H[43]), .A2(n148), .B0(n663), 
        .B1(n122), .Y(MULi_1_mult_15_n84) );
  OAI32X4 U546 ( .A0(SR_to_MUL[48]), .A1(TEMP_H[50]), .A2(n149), .B0(n281), 
        .B1(n288), .Y(MULi_0_mult_15_n85) );
  OAI32X4 U547 ( .A0(SR_to_MUL[48]), .A1(TEMP_H[51]), .A2(n149), .B0(n279), 
        .B1(n123), .Y(MULi_0_mult_15_n84) );
  OAI22X2 U548 ( .A0(n78), .A1(n459), .B0(n462), .B1(n463), .Y(
        MULi_4_mult_15_n77) );
  OAI32X4 U549 ( .A0(n460), .A1(n105), .A2(n78), .B0(n462), .B1(n460), .Y(
        MULi_4_mult_15_n54) );
  OAI22X2 U550 ( .A0(n78), .A1(n457), .B0(n462), .B1(n458), .Y(
        MULi_4_mult_15_n75) );
  OAI22X2 U551 ( .A0(n78), .A1(n456), .B0(n462), .B1(n457), .Y(
        MULi_4_mult_15_n74) );
  INVX6 U552 ( .A(n170), .Y(n462) );
  OAI22X2 U553 ( .A0(n79), .A1(n394), .B0(n398), .B1(n395), .Y(
        MULi_5_mult_15_n76) );
  OAI32X4 U554 ( .A0(n396), .A1(n107), .A2(n79), .B0(n398), .B1(n396), .Y(
        MULi_5_mult_15_n54) );
  OAI22X2 U555 ( .A0(n79), .A1(n393), .B0(n398), .B1(n394), .Y(
        MULi_5_mult_15_n75) );
  OAI22X2 U556 ( .A0(n79), .A1(n392), .B0(n398), .B1(n393), .Y(
        MULi_5_mult_15_n74) );
  INVX6 U557 ( .A(n172), .Y(n398) );
  OAI22X2 U558 ( .A0(n74), .A1(n523), .B0(n526), .B1(n527), .Y(
        MULi_3_mult_15_n77) );
  OAI22X2 U559 ( .A0(n74), .A1(n522), .B0(n526), .B1(n523), .Y(
        MULi_3_mult_15_n76) );
  OAI32X4 U560 ( .A0(n524), .A1(n104), .A2(n74), .B0(n526), .B1(n524), .Y(
        MULi_3_mult_15_n54) );
  OAI22X2 U561 ( .A0(n74), .A1(n521), .B0(n526), .B1(n522), .Y(
        MULi_3_mult_15_n75) );
  OAI22X2 U562 ( .A0(n74), .A1(n520), .B0(n526), .B1(n521), .Y(
        MULi_3_mult_15_n74) );
  INVX6 U563 ( .A(n171), .Y(n526) );
  OAI22X2 U564 ( .A0(n80), .A1(n331), .B0(n334), .B1(n335), .Y(
        MULi_6_mult_15_n77) );
  OAI22X2 U565 ( .A0(n80), .A1(n330), .B0(n334), .B1(n331), .Y(
        MULi_6_mult_15_n76) );
  OAI32X4 U566 ( .A0(n332), .A1(n109), .A2(n80), .B0(n334), .B1(n332), .Y(
        MULi_6_mult_15_n54) );
  OAI22X2 U567 ( .A0(n80), .A1(n329), .B0(n334), .B1(n330), .Y(
        MULi_6_mult_15_n75) );
  OAI22X2 U568 ( .A0(n80), .A1(n328), .B0(n334), .B1(n329), .Y(
        MULi_6_mult_15_n74) );
  INVX6 U569 ( .A(n326), .Y(n334) );
  OAI22X2 U570 ( .A0(n77), .A1(n587), .B0(n590), .B1(n591), .Y(
        MULi_2_mult_15_n77) );
  OAI32X4 U571 ( .A0(n588), .A1(n106), .A2(n77), .B0(n590), .B1(n588), .Y(
        MULi_2_mult_15_n54) );
  OAI22X2 U572 ( .A0(n77), .A1(n585), .B0(n590), .B1(n586), .Y(
        MULi_2_mult_15_n75) );
  OAI22X2 U573 ( .A0(n77), .A1(n584), .B0(n590), .B1(n585), .Y(
        MULi_2_mult_15_n74) );
  INVX6 U574 ( .A(n173), .Y(n590) );
  OAI22X2 U575 ( .A0(n76), .A1(n267), .B0(n270), .B1(n271), .Y(
        MULi_0_mult_15_n77) );
  OAI22X2 U576 ( .A0(n76), .A1(n266), .B0(n270), .B1(n267), .Y(
        MULi_0_mult_15_n76) );
  OAI32X4 U577 ( .A0(n268), .A1(n110), .A2(n76), .B0(n270), .B1(n268), .Y(
        MULi_0_mult_15_n54) );
  OAI22X2 U578 ( .A0(n76), .A1(n265), .B0(n270), .B1(n266), .Y(
        MULi_0_mult_15_n75) );
  OAI22X2 U579 ( .A0(n76), .A1(n264), .B0(n270), .B1(n265), .Y(
        MULi_0_mult_15_n74) );
  INVX6 U580 ( .A(n174), .Y(n270) );
  OAI32X4 U581 ( .A0(n652), .A1(n108), .A2(n75), .B0(n654), .B1(n652), .Y(
        MULi_1_mult_15_n54) );
  OAI22X2 U582 ( .A0(n75), .A1(n649), .B0(n654), .B1(n650), .Y(
        MULi_1_mult_15_n75) );
  OAI22X2 U583 ( .A0(n75), .A1(n648), .B0(n654), .B1(n649), .Y(
        MULi_1_mult_15_n74) );
  INVX6 U584 ( .A(n175), .Y(n654) );
  AOI22X4 U585 ( .A0(n546), .A1(n538), .B0(TEMP_H[26]), .B1(n512), .Y(n511) );
  AOI22X4 U586 ( .A0(n547), .A1(n538), .B0(TEMP_H[26]), .B1(n524), .Y(n523) );
  AOI22X4 U587 ( .A0(n546), .A1(n534), .B0(TEMP_H[28]), .B1(n512), .Y(n509) );
  AOI22X4 U588 ( .A0(n547), .A1(n534), .B0(TEMP_H[28]), .B1(n524), .Y(n521) );
  AOI22X4 U589 ( .A0(n482), .A1(n470), .B0(TEMP_H[20]), .B1(n448), .Y(n445) );
  AOI22X4 U590 ( .A0(n483), .A1(n470), .B0(TEMP_H[20]), .B1(n460), .Y(n457) );
  AOI22X4 U591 ( .A0(n610), .A1(n602), .B0(TEMP_H[34]), .B1(n576), .Y(n575) );
  AOI22X4 U592 ( .A0(n611), .A1(n602), .B0(TEMP_H[34]), .B1(n588), .Y(n587) );
  AOI22X4 U593 ( .A0(n482), .A1(n474), .B0(TEMP_H[18]), .B1(n448), .Y(n447) );
  AOI22X4 U594 ( .A0(n483), .A1(n474), .B0(TEMP_H[18]), .B1(n460), .Y(n459) );
  AOI22X4 U595 ( .A0(n610), .A1(n598), .B0(TEMP_H[36]), .B1(n576), .Y(n573) );
  AOI22X4 U596 ( .A0(n611), .A1(n598), .B0(TEMP_H[36]), .B1(n588), .Y(n585) );
  AOI22X4 U597 ( .A0(n418), .A1(n406), .B0(TEMP_H[12]), .B1(n384), .Y(n381) );
  AOI22X4 U598 ( .A0(n419), .A1(n406), .B0(TEMP_H[12]), .B1(n396), .Y(n393) );
  AOI22X4 U599 ( .A0(n674), .A1(n666), .B0(TEMP_H[42]), .B1(n640), .Y(n639) );
  AOI22X4 U600 ( .A0(n675), .A1(n666), .B0(TEMP_H[42]), .B1(n652), .Y(n651) );
  AOI22X4 U601 ( .A0(n418), .A1(n410), .B0(TEMP_H[10]), .B1(n384), .Y(n383) );
  AOI22X4 U602 ( .A0(n419), .A1(n410), .B0(TEMP_H[10]), .B1(n396), .Y(n395) );
  AOI22X4 U603 ( .A0(n674), .A1(n662), .B0(TEMP_H[44]), .B1(n640), .Y(n637) );
  AOI22X4 U604 ( .A0(n675), .A1(n662), .B0(TEMP_H[44]), .B1(n652), .Y(n649) );
  AOI22X4 U605 ( .A0(n354), .A1(n344), .B0(TEMP_H[3]), .B1(n320), .Y(n318) );
  AOI22X4 U606 ( .A0(n355), .A1(n344), .B0(TEMP_H[3]), .B1(n332), .Y(n330) );
  AOI22X4 U607 ( .A0(n290), .A1(n282), .B0(TEMP_H[50]), .B1(n256), .Y(n255) );
  AOI22X4 U608 ( .A0(n291), .A1(n282), .B0(TEMP_H[50]), .B1(n268), .Y(n267) );
  AOI22X4 U609 ( .A0(n354), .A1(n346), .B0(TEMP_H[2]), .B1(n320), .Y(n319) );
  AOI22X4 U610 ( .A0(n355), .A1(n346), .B0(TEMP_H[2]), .B1(n332), .Y(n331) );
  AOI22X4 U611 ( .A0(n290), .A1(n278), .B0(TEMP_H[52]), .B1(n256), .Y(n253) );
  AOI22X4 U612 ( .A0(n291), .A1(n278), .B0(TEMP_H[52]), .B1(n268), .Y(n265) );
  AOI22X4 U613 ( .A0(n355), .A1(n342), .B0(TEMP_H[4]), .B1(n332), .Y(n329) );
  OAI32X4 U614 ( .A0(n111), .A1(TEMP_H[30]), .A2(n152), .B0(n529), .B1(n118), 
        .Y(MULi_3_mult_15_n81) );
  AOI22X4 U615 ( .A0(TEMP_H[30]), .A1(n512), .B0(n546), .B1(n530), .Y(n507) );
  OAI32X4 U616 ( .A0(n113), .A1(TEMP_H[22]), .A2(n154), .B0(n465), .B1(n117), 
        .Y(MULi_4_mult_15_n81) );
  AOI22X4 U617 ( .A0(TEMP_H[22]), .A1(n448), .B0(n482), .B1(n466), .Y(n443) );
  OAI32X4 U618 ( .A0(n112), .A1(TEMP_H[38]), .A2(n153), .B0(n593), .B1(n120), 
        .Y(MULi_2_mult_15_n81) );
  AOI22X4 U619 ( .A0(TEMP_H[38]), .A1(n576), .B0(n610), .B1(n594), .Y(n571) );
  OAI32X4 U620 ( .A0(n115), .A1(TEMP_H[14]), .A2(n151), .B0(n401), .B1(n119), 
        .Y(MULi_5_mult_15_n81) );
  AOI22X4 U621 ( .A0(TEMP_H[14]), .A1(n384), .B0(n418), .B1(n402), .Y(n379) );
  OAI32X4 U622 ( .A0(n114), .A1(TEMP_H[46]), .A2(n148), .B0(n657), .B1(n122), 
        .Y(MULi_1_mult_15_n81) );
  AOI22X4 U623 ( .A0(TEMP_H[46]), .A1(n640), .B0(n674), .B1(n658), .Y(n635) );
  OAI32X4 U624 ( .A0(n103), .A1(TEMP_H[6]), .A2(n150), .B0(n337), .B1(n121), 
        .Y(MULi_6_mult_15_n81) );
  AOI22X4 U625 ( .A0(TEMP_H[6]), .A1(n320), .B0(n354), .B1(n338), .Y(n315) );
  OAI32X4 U626 ( .A0(n116), .A1(TEMP_H[54]), .A2(n149), .B0(n273), .B1(n123), 
        .Y(MULi_0_mult_15_n81) );
  AOI22X4 U627 ( .A0(TEMP_H[54]), .A1(n256), .B0(n290), .B1(n274), .Y(n251) );
  AOI22X4 U628 ( .A0(n547), .A1(n536), .B0(TEMP_H[27]), .B1(n524), .Y(n522) );
  AOI22X4 U629 ( .A0(n611), .A1(n600), .B0(TEMP_H[35]), .B1(n588), .Y(n586) );
  AOI22X4 U630 ( .A0(n483), .A1(n472), .B0(TEMP_H[19]), .B1(n460), .Y(n458) );
  AOI22X4 U631 ( .A0(n675), .A1(n664), .B0(TEMP_H[43]), .B1(n652), .Y(n650) );
  AOI22X4 U632 ( .A0(n419), .A1(n408), .B0(TEMP_H[11]), .B1(n396), .Y(n394) );
  AOI22X4 U633 ( .A0(n291), .A1(n280), .B0(TEMP_H[51]), .B1(n268), .Y(n266) );
  AOI22X4 U634 ( .A0(TEMP_H[29]), .A1(n512), .B0(n546), .B1(n532), .Y(n508) );
  OAI22X4 U635 ( .A0(n524), .A1(n532), .B0(TEMP_H[29]), .B1(n547), .Y(n520) );
  OAI32X4 U636 ( .A0(n111), .A1(TEMP_H[29]), .A2(n152), .B0(n531), .B1(n118), 
        .Y(MULi_3_mult_15_n82) );
  AOI22X4 U637 ( .A0(TEMP_H[37]), .A1(n576), .B0(n610), .B1(n596), .Y(n572) );
  OAI22X4 U638 ( .A0(n588), .A1(n596), .B0(TEMP_H[37]), .B1(n611), .Y(n584) );
  OAI32X4 U639 ( .A0(n112), .A1(TEMP_H[37]), .A2(n153), .B0(n595), .B1(n120), 
        .Y(MULi_2_mult_15_n82) );
  AOI22X4 U640 ( .A0(TEMP_H[21]), .A1(n448), .B0(n482), .B1(n468), .Y(n444) );
  OAI22X4 U641 ( .A0(n460), .A1(n468), .B0(TEMP_H[21]), .B1(n483), .Y(n456) );
  OAI32X4 U642 ( .A0(n113), .A1(TEMP_H[21]), .A2(n154), .B0(n467), .B1(n117), 
        .Y(MULi_4_mult_15_n82) );
  AOI22X4 U643 ( .A0(TEMP_H[45]), .A1(n640), .B0(n674), .B1(n660), .Y(n636) );
  OAI22X4 U644 ( .A0(n652), .A1(n660), .B0(TEMP_H[45]), .B1(n675), .Y(n648) );
  OAI32X4 U645 ( .A0(n114), .A1(TEMP_H[45]), .A2(n148), .B0(n659), .B1(n122), 
        .Y(MULi_1_mult_15_n82) );
  AOI22X4 U646 ( .A0(TEMP_H[13]), .A1(n384), .B0(n418), .B1(n404), .Y(n380) );
  OAI22X4 U647 ( .A0(n396), .A1(n404), .B0(TEMP_H[13]), .B1(n419), .Y(n392) );
  OAI32X4 U648 ( .A0(n115), .A1(TEMP_H[13]), .A2(n151), .B0(n403), .B1(n119), 
        .Y(MULi_5_mult_15_n82) );
  AOI22X4 U649 ( .A0(TEMP_H[53]), .A1(n256), .B0(n290), .B1(n276), .Y(n252) );
  OAI22X4 U650 ( .A0(n268), .A1(n276), .B0(TEMP_H[53]), .B1(n291), .Y(n264) );
  OAI32X4 U651 ( .A0(n116), .A1(TEMP_H[53]), .A2(n149), .B0(n275), .B1(n123), 
        .Y(MULi_0_mult_15_n82) );
  AOI22X4 U652 ( .A0(TEMP_H[5]), .A1(n320), .B0(n354), .B1(n340), .Y(n316) );
  OAI22X4 U653 ( .A0(n332), .A1(n340), .B0(TEMP_H[5]), .B1(n355), .Y(n328) );
  OAI32X4 U654 ( .A0(n103), .A1(TEMP_H[5]), .A2(n150), .B0(n339), .B1(n121), 
        .Y(MULi_6_mult_15_n82) );
  BUFX10 U655 ( .A(SR_to_MUL[29]), .Y(n546) );
  BUFX10 U656 ( .A(SR_to_MUL[21]), .Y(n482) );
  BUFX10 U657 ( .A(SR_to_MUL[37]), .Y(n610) );
  BUFX10 U658 ( .A(SR_to_MUL[13]), .Y(n418) );
  BUFX10 U659 ( .A(SR_to_MUL[45]), .Y(n674) );
  BUFX10 U660 ( .A(SR_to_MUL[53]), .Y(n290) );
  BUFX10 U661 ( .A(SR_to_MUL[5]), .Y(n354) );
  BUFX10 U662 ( .A(SR_to_MUL[19]), .Y(n483) );
  BUFX10 U663 ( .A(SR_to_MUL[27]), .Y(n547) );
  BUFX10 U664 ( .A(SR_to_MUL[11]), .Y(n419) );
  BUFX10 U665 ( .A(SR_to_MUL[35]), .Y(n611) );
  BUFX10 U666 ( .A(SR_to_MUL[43]), .Y(n675) );
  BUFX10 U667 ( .A(SR_to_MUL[51]), .Y(n291) );
  OAI32X4 U668 ( .A0(n512), .A1(n104), .A2(n551), .B0(n552), .B1(n512), .Y(
        MULi_3_mult_15_n53) );
  OAI32X4 U669 ( .A0(n576), .A1(n106), .A2(n615), .B0(n616), .B1(n576), .Y(
        MULi_2_mult_15_n53) );
  OAI32X4 U670 ( .A0(n448), .A1(n105), .A2(n487), .B0(n488), .B1(n448), .Y(
        MULi_4_mult_15_n53) );
  OAI32X4 U671 ( .A0(n640), .A1(n108), .A2(n679), .B0(n680), .B1(n640), .Y(
        MULi_1_mult_15_n53) );
  OAI32X4 U672 ( .A0(n384), .A1(n107), .A2(n423), .B0(n424), .B1(n384), .Y(
        MULi_5_mult_15_n53) );
  OAI32X4 U673 ( .A0(n256), .A1(n110), .A2(n295), .B0(n296), .B1(n256), .Y(
        MULi_0_mult_15_n53) );
  OAI32X4 U674 ( .A0(n320), .A1(n109), .A2(n359), .B0(n360), .B1(n320), .Y(
        MULi_6_mult_15_n53) );
  AOI22X4 U675 ( .A0(n354), .A1(n342), .B0(TEMP_H[4]), .B1(n320), .Y(n317) );
  AOI22X4 U676 ( .A0(TEMP_H[5]), .A1(n309), .B0(n353), .B1(n340), .Y(n305) );
  AOI22X4 U677 ( .A0(TEMP_H[13]), .A1(n373), .B0(n417), .B1(n404), .Y(n369) );
  AOI22X4 U678 ( .A0(TEMP_H[21]), .A1(n437), .B0(n481), .B1(n468), .Y(n433) );
  AOI22X4 U679 ( .A0(TEMP_H[37]), .A1(n565), .B0(n609), .B1(n596), .Y(n561) );
  AOI22X4 U680 ( .A0(TEMP_H[53]), .A1(n245), .B0(n289), .B1(n276), .Y(n241) );
  AOI22X4 U681 ( .A0(TEMP_H[45]), .A1(n629), .B0(n673), .B1(n660), .Y(n625) );
  AOI22X4 U682 ( .A0(TEMP_H[29]), .A1(n501), .B0(n545), .B1(n532), .Y(n497) );
  AOI22X4 U683 ( .A0(TEMP_H[7]), .A1(n320), .B0(n354), .B1(n336), .Y(n314) );
  AOI22X4 U684 ( .A0(n418), .A1(n408), .B0(TEMP_H[11]), .B1(n384), .Y(n382) );
  AOI22X4 U685 ( .A0(n482), .A1(n472), .B0(TEMP_H[19]), .B1(n448), .Y(n446) );
  AOI22X4 U686 ( .A0(n610), .A1(n600), .B0(TEMP_H[35]), .B1(n576), .Y(n574) );
  AOI22X4 U687 ( .A0(n290), .A1(n280), .B0(TEMP_H[51]), .B1(n256), .Y(n254) );
  AOI22X4 U688 ( .A0(n674), .A1(n664), .B0(TEMP_H[43]), .B1(n640), .Y(n638) );
  AOI22X4 U689 ( .A0(n546), .A1(n536), .B0(TEMP_H[27]), .B1(n512), .Y(n510) );
  AOI22X4 U690 ( .A0(TEMP_H[6]), .A1(n355), .B0(n332), .B1(n338), .Y(n300) );
  AOI22X4 U691 ( .A0(TEMP_H[14]), .A1(n419), .B0(n396), .B1(n402), .Y(n364) );
  AOI22X4 U692 ( .A0(TEMP_H[22]), .A1(n483), .B0(n460), .B1(n466), .Y(n428) );
  AOI22X4 U693 ( .A0(TEMP_H[38]), .A1(n611), .B0(n588), .B1(n594), .Y(n556) );
  AOI22X4 U694 ( .A0(TEMP_H[54]), .A1(n291), .B0(n268), .B1(n274), .Y(n236) );
  AOI22X4 U695 ( .A0(TEMP_H[46]), .A1(n675), .B0(n652), .B1(n658), .Y(n620) );
  AOI22X4 U696 ( .A0(TEMP_H[30]), .A1(n547), .B0(n524), .B1(n530), .Y(n492) );
  OAI22X4 U697 ( .A0(n357), .A1(n303), .B0(n358), .B1(n304), .Y(
        MULi_6_mult_15_n15) );
  OAI22X4 U698 ( .A0(n421), .A1(n367), .B0(n422), .B1(n368), .Y(
        MULi_5_mult_15_n15) );
  OAI22X4 U699 ( .A0(n485), .A1(n431), .B0(n486), .B1(n432), .Y(
        MULi_4_mult_15_n15) );
  OAI22X4 U700 ( .A0(n613), .A1(n559), .B0(n614), .B1(n560), .Y(
        MULi_2_mult_15_n15) );
  OAI22X4 U701 ( .A0(n293), .A1(n239), .B0(n294), .B1(n240), .Y(
        MULi_0_mult_15_n15) );
  OAI22X4 U702 ( .A0(n677), .A1(n623), .B0(n678), .B1(n624), .Y(
        MULi_1_mult_15_n15) );
  OAI22X4 U703 ( .A0(n549), .A1(n495), .B0(n550), .B1(n496), .Y(
        MULi_3_mult_15_n15) );
  OAI22X4 U704 ( .A0(n423), .A1(n378), .B0(n424), .B1(n379), .Y(
        MULi_5_mult_15_n21) );
  OAI22X4 U705 ( .A0(n487), .A1(n442), .B0(n488), .B1(n443), .Y(
        MULi_4_mult_15_n21) );
  OAI22X4 U706 ( .A0(n615), .A1(n570), .B0(n616), .B1(n571), .Y(
        MULi_2_mult_15_n21) );
  OAI22X4 U707 ( .A0(n295), .A1(n250), .B0(n296), .B1(n251), .Y(
        MULi_0_mult_15_n21) );
  OAI22X4 U708 ( .A0(n679), .A1(n634), .B0(n680), .B1(n635), .Y(
        MULi_1_mult_15_n21) );
  OAI22X4 U709 ( .A0(n551), .A1(n506), .B0(n552), .B1(n507), .Y(
        MULi_3_mult_15_n21) );
  INVX2 U710 ( .A(n336), .Y(n180) );
  INVX2 U711 ( .A(TEMP_H[7]), .Y(n181) );
  XNOR2X2 U712 ( .A(n302), .B(n301), .Y(MULi_6_mult_15_n35) );
  INVX2 U713 ( .A(n400), .Y(n186) );
  INVX2 U714 ( .A(TEMP_H[15]), .Y(n187) );
  XNOR2X2 U715 ( .A(n366), .B(n365), .Y(MULi_5_mult_15_n35) );
  INVX2 U716 ( .A(n464), .Y(n192) );
  INVX2 U717 ( .A(TEMP_H[23]), .Y(n193) );
  XNOR2X2 U718 ( .A(n430), .B(n429), .Y(MULi_4_mult_15_n35) );
  INVX2 U719 ( .A(n592), .Y(n198) );
  INVX2 U720 ( .A(TEMP_H[39]), .Y(n199) );
  XNOR2X2 U721 ( .A(n558), .B(n557), .Y(MULi_2_mult_15_n35) );
  INVX2 U722 ( .A(n272), .Y(n204) );
  INVX2 U723 ( .A(TEMP_H[55]), .Y(n205) );
  XNOR2X2 U724 ( .A(n238), .B(n237), .Y(MULi_0_mult_15_n35) );
  INVX2 U725 ( .A(n656), .Y(n210) );
  INVX2 U726 ( .A(TEMP_H[47]), .Y(n211) );
  XNOR2X2 U727 ( .A(n622), .B(n621), .Y(MULi_1_mult_15_n35) );
  INVX2 U728 ( .A(n528), .Y(n216) );
  INVX2 U729 ( .A(TEMP_H[31]), .Y(n217) );
  XNOR2X2 U730 ( .A(n494), .B(n493), .Y(MULi_3_mult_15_n35) );
  AOI22X2 U731 ( .A0(TEMP_H[52]), .A1(n245), .B0(n289), .B1(n278), .Y(n242) );
  AOI22X2 U732 ( .A0(n290), .A1(n283), .B0(TEMP_H[49]), .B1(n256), .Y(n259) );
  AOI22X1 U733 ( .A0(n292), .A1(n282), .B0(TEMP_H[50]), .B1(n149), .Y(n284) );
  AOI22X2 U734 ( .A0(n292), .A1(n283), .B0(TEMP_H[49]), .B1(n149), .Y(n285) );
  AOI22X2 U735 ( .A0(n291), .A1(TEMP_H[55]), .B0(n272), .B1(n268), .Y(n261) );
  OAI21X1 U736 ( .A0(n263), .A1(n174), .B0(n261), .Y(MULi_0_mult_15_n72) );
  AOI22X2 U737 ( .A0(TEMP_H[49]), .A1(n245), .B0(n289), .B1(n283), .Y(n248) );
  AOI22X2 U738 ( .A0(TEMP_H[50]), .A1(n245), .B0(n289), .B1(n282), .Y(n244) );
  AOI22X2 U739 ( .A0(TEMP_H[51]), .A1(n245), .B0(n289), .B1(n280), .Y(n243) );
  OAI22X1 U740 ( .A0(n293), .A1(n240), .B0(n294), .B1(n241), .Y(
        MULi_0_mult_15_n57) );
  OAI22X1 U741 ( .A0(n293), .A1(n241), .B0(n294), .B1(n242), .Y(
        MULi_0_mult_15_n58) );
  OAI22X1 U742 ( .A0(n295), .A1(n259), .B0(n296), .B1(n257), .Y(
        MULi_0_mult_15_n70) );
  OAI22X1 U743 ( .A0(n288), .A1(n284), .B0(n286), .B1(n285), .Y(
        MULi_0_mult_15_n86) );
  AOI21X1 U744 ( .A0(SR_to_MUL[48]), .A1(TEMP_H[48]), .B0(n149), .Y(
        MULi_0_mult_15_n55) );
  OAI22X1 U745 ( .A0(TEMP_H[48]), .A1(n286), .B0(n288), .B1(n285), .Y(
        MULi_0_mult_15_n87) );
  OAI22X1 U746 ( .A0(n293), .A1(n248), .B0(n294), .B1(n246), .Y(
        MULi_0_mult_15_n62) );
  OAI22X1 U747 ( .A0(n295), .A1(n255), .B0(n296), .B1(n259), .Y(
        MULi_0_mult_15_n69) );
  OAI22X1 U748 ( .A0(n295), .A1(n254), .B0(n296), .B1(n255), .Y(
        MULi_0_mult_15_n68) );
  OAI22X1 U749 ( .A0(n293), .A1(n244), .B0(n248), .B1(n294), .Y(
        MULi_0_mult_15_n61) );
  OAI22X1 U750 ( .A0(n295), .A1(n253), .B0(n296), .B1(n254), .Y(
        MULi_0_mult_15_n67) );
  OAI22X1 U751 ( .A0(n293), .A1(n243), .B0(n294), .B1(n244), .Y(
        MULi_0_mult_15_n60) );
  OAI22X1 U752 ( .A0(n295), .A1(n252), .B0(n296), .B1(n253), .Y(
        MULi_0_mult_15_n66) );
  OAI22X1 U753 ( .A0(n295), .A1(n251), .B0(n296), .B1(n252), .Y(
        MULi_0_mult_15_n65) );
  OAI22X1 U754 ( .A0(n293), .A1(n242), .B0(n294), .B1(n243), .Y(
        MULi_0_mult_15_n59) );
  INVX4 U755 ( .A(n76), .Y(n263) );
  AOI22X2 U756 ( .A0(n354), .A1(n347), .B0(TEMP_H[1]), .B1(n320), .Y(n323) );
  AOI22X2 U757 ( .A0(n355), .A1(TEMP_H[7]), .B0(n336), .B1(n332), .Y(n325) );
  AOI22X2 U758 ( .A0(TEMP_H[1]), .A1(n309), .B0(n353), .B1(n347), .Y(n312) );
  AOI22X2 U759 ( .A0(TEMP_H[2]), .A1(n309), .B0(n353), .B1(n346), .Y(n308) );
  AOI22X2 U760 ( .A0(TEMP_H[3]), .A1(n309), .B0(n353), .B1(n344), .Y(n307) );
  OAI22X1 U761 ( .A0(n357), .A1(n304), .B0(n358), .B1(n305), .Y(
        MULi_6_mult_15_n57) );
  OAI22X1 U762 ( .A0(n357), .A1(n305), .B0(n358), .B1(n155), .Y(
        MULi_6_mult_15_n58) );
  OAI22X1 U763 ( .A0(n359), .A1(n323), .B0(n360), .B1(n321), .Y(
        MULi_6_mult_15_n70) );
  AOI22X1 U764 ( .A0(n356), .A1(n346), .B0(TEMP_H[2]), .B1(n150), .Y(n348) );
  AOI22X2 U765 ( .A0(n356), .A1(n347), .B0(TEMP_H[1]), .B1(n150), .Y(n349) );
  OAI22X1 U766 ( .A0(n352), .A1(n348), .B0(n350), .B1(n349), .Y(
        MULi_6_mult_15_n86) );
  AOI21X1 U767 ( .A0(SR_to_MUL[0]), .A1(TEMP_H[0]), .B0(n150), .Y(
        MULi_6_mult_15_n55) );
  OAI22X1 U768 ( .A0(TEMP_H[0]), .A1(n350), .B0(n352), .B1(n349), .Y(
        MULi_6_mult_15_n87) );
  ADDFX1 U769 ( .A(MULi_6_mult_15_n19), .B(MULi_6_mult_15_n18), .CI(
        MULi_6_mult_15_n4), .CO(MULi_6_mult_15_n3), .S(MUL_to_PIPE1[12]) );
  ADDFX1 U770 ( .A(MULi_6_mult_15_n17), .B(MULi_6_mult_15_n16), .CI(
        MULi_6_mult_15_n3), .CO(MULi_6_mult_15_n2), .S(MUL_to_PIPE1[13]) );
  ADDFX1 U771 ( .A(MULi_6_mult_15_n15), .B(MULi_6_mult_15_n56), .CI(
        MULi_6_mult_15_n2), .CO(MULi_6_mult_15_n1), .S(MUL_to_PIPE1[14]) );
  OAI21X1 U772 ( .A0(n327), .A1(n176), .B0(n325), .Y(MULi_6_mult_15_n72) );
  OAI22X1 U773 ( .A0(n357), .A1(n312), .B0(n358), .B1(n310), .Y(
        MULi_6_mult_15_n62) );
  OAI22X1 U774 ( .A0(n359), .A1(n319), .B0(n360), .B1(n323), .Y(
        MULi_6_mult_15_n69) );
  OAI22X1 U775 ( .A0(n359), .A1(n318), .B0(n360), .B1(n319), .Y(
        MULi_6_mult_15_n68) );
  OAI22X1 U776 ( .A0(n357), .A1(n308), .B0(n312), .B1(n358), .Y(
        MULi_6_mult_15_n61) );
  OAI22X1 U777 ( .A0(n359), .A1(n317), .B0(n360), .B1(n318), .Y(
        MULi_6_mult_15_n67) );
  OAI22X1 U778 ( .A0(n357), .A1(n307), .B0(n358), .B1(n308), .Y(
        MULi_6_mult_15_n60) );
  OAI22X1 U779 ( .A0(n359), .A1(n315), .B0(n360), .B1(n316), .Y(
        MULi_6_mult_15_n65) );
  OAI22X1 U780 ( .A0(n357), .A1(n306), .B0(n358), .B1(n307), .Y(
        MULi_6_mult_15_n59) );
  AOI22X2 U781 ( .A0(TEMP_H[12]), .A1(n373), .B0(n417), .B1(n406), .Y(n370) );
  AOI22X2 U782 ( .A0(n418), .A1(n411), .B0(TEMP_H[9]), .B1(n384), .Y(n387) );
  AOI22X1 U783 ( .A0(n420), .A1(n410), .B0(TEMP_H[10]), .B1(n151), .Y(n412) );
  AOI22X2 U784 ( .A0(n420), .A1(n411), .B0(TEMP_H[9]), .B1(n151), .Y(n413) );
  AOI22X2 U785 ( .A0(n419), .A1(TEMP_H[15]), .B0(n400), .B1(n396), .Y(n389) );
  OAI21X1 U786 ( .A0(n391), .A1(n172), .B0(n389), .Y(MULi_5_mult_15_n72) );
  AOI22X2 U787 ( .A0(TEMP_H[9]), .A1(n373), .B0(n417), .B1(n411), .Y(n376) );
  AOI22X2 U788 ( .A0(TEMP_H[10]), .A1(n373), .B0(n417), .B1(n410), .Y(n372) );
  AOI22X2 U789 ( .A0(TEMP_H[11]), .A1(n373), .B0(n417), .B1(n408), .Y(n371) );
  OAI22X1 U790 ( .A0(n421), .A1(n368), .B0(n422), .B1(n369), .Y(
        MULi_5_mult_15_n57) );
  OAI22X1 U791 ( .A0(n421), .A1(n369), .B0(n422), .B1(n370), .Y(
        MULi_5_mult_15_n58) );
  OAI22X1 U792 ( .A0(n423), .A1(n387), .B0(n424), .B1(n385), .Y(
        MULi_5_mult_15_n70) );
  OAI22X1 U793 ( .A0(n416), .A1(n412), .B0(n414), .B1(n413), .Y(
        MULi_5_mult_15_n86) );
  AOI21X1 U794 ( .A0(SR_to_MUL[8]), .A1(TEMP_H[8]), .B0(n151), .Y(
        MULi_5_mult_15_n55) );
  OAI22X1 U795 ( .A0(TEMP_H[8]), .A1(n414), .B0(n416), .B1(n413), .Y(
        MULi_5_mult_15_n87) );
  ADDFX1 U796 ( .A(MULi_5_mult_15_n19), .B(MULi_5_mult_15_n18), .CI(
        MULi_5_mult_15_n4), .CO(MULi_5_mult_15_n3), .S(MUL_to_PIPE1[28]) );
  ADDFX1 U797 ( .A(MULi_5_mult_15_n17), .B(MULi_5_mult_15_n16), .CI(
        MULi_5_mult_15_n3), .CO(MULi_5_mult_15_n2), .S(MUL_to_PIPE1[29]) );
  ADDFX1 U798 ( .A(MULi_5_mult_15_n15), .B(MULi_5_mult_15_n56), .CI(
        MULi_5_mult_15_n2), .CO(MULi_5_mult_15_n1), .S(MUL_to_PIPE1[30]) );
  OAI22X1 U799 ( .A0(n421), .A1(n376), .B0(n422), .B1(n374), .Y(
        MULi_5_mult_15_n62) );
  OAI22X1 U800 ( .A0(n423), .A1(n383), .B0(n424), .B1(n387), .Y(
        MULi_5_mult_15_n69) );
  OAI22X1 U801 ( .A0(n423), .A1(n382), .B0(n424), .B1(n383), .Y(
        MULi_5_mult_15_n68) );
  OAI22X1 U802 ( .A0(n421), .A1(n372), .B0(n376), .B1(n422), .Y(
        MULi_5_mult_15_n61) );
  OAI22X1 U803 ( .A0(n423), .A1(n381), .B0(n424), .B1(n382), .Y(
        MULi_5_mult_15_n67) );
  OAI22X1 U804 ( .A0(n421), .A1(n371), .B0(n422), .B1(n372), .Y(
        MULi_5_mult_15_n60) );
  OAI22X1 U805 ( .A0(n423), .A1(n380), .B0(n424), .B1(n381), .Y(
        MULi_5_mult_15_n66) );
  OAI22X1 U806 ( .A0(n423), .A1(n379), .B0(n424), .B1(n380), .Y(
        MULi_5_mult_15_n65) );
  OAI22X1 U807 ( .A0(n421), .A1(n370), .B0(n422), .B1(n371), .Y(
        MULi_5_mult_15_n59) );
  INVX4 U808 ( .A(n79), .Y(n391) );
  AOI22X2 U809 ( .A0(TEMP_H[20]), .A1(n437), .B0(n481), .B1(n470), .Y(n434) );
  AOI22X2 U810 ( .A0(n482), .A1(n475), .B0(TEMP_H[17]), .B1(n448), .Y(n451) );
  AOI22X1 U811 ( .A0(n484), .A1(n474), .B0(TEMP_H[18]), .B1(n154), .Y(n476) );
  AOI22X2 U812 ( .A0(n484), .A1(n475), .B0(TEMP_H[17]), .B1(n154), .Y(n477) );
  AOI22X2 U813 ( .A0(n483), .A1(TEMP_H[23]), .B0(n464), .B1(n460), .Y(n453) );
  OAI21X1 U814 ( .A0(n455), .A1(n170), .B0(n453), .Y(MULi_4_mult_15_n72) );
  AOI22X2 U815 ( .A0(TEMP_H[17]), .A1(n437), .B0(n481), .B1(n475), .Y(n440) );
  AOI22X2 U816 ( .A0(TEMP_H[18]), .A1(n437), .B0(n481), .B1(n474), .Y(n436) );
  AOI22X2 U817 ( .A0(TEMP_H[19]), .A1(n437), .B0(n481), .B1(n472), .Y(n435) );
  OAI22X1 U818 ( .A0(n485), .A1(n432), .B0(n486), .B1(n433), .Y(
        MULi_4_mult_15_n57) );
  OAI22X1 U819 ( .A0(n485), .A1(n433), .B0(n486), .B1(n434), .Y(
        MULi_4_mult_15_n58) );
  OAI22X1 U820 ( .A0(n487), .A1(n451), .B0(n488), .B1(n449), .Y(
        MULi_4_mult_15_n70) );
  OAI22X1 U821 ( .A0(n480), .A1(n476), .B0(n478), .B1(n477), .Y(
        MULi_4_mult_15_n86) );
  AOI21X1 U822 ( .A0(SR_to_MUL[16]), .A1(TEMP_H[16]), .B0(n154), .Y(
        MULi_4_mult_15_n55) );
  OAI22X1 U823 ( .A0(TEMP_H[16]), .A1(n478), .B0(n480), .B1(n477), .Y(
        MULi_4_mult_15_n87) );
  OAI22X1 U824 ( .A0(n485), .A1(n440), .B0(n486), .B1(n438), .Y(
        MULi_4_mult_15_n62) );
  OAI22X1 U825 ( .A0(n487), .A1(n447), .B0(n488), .B1(n451), .Y(
        MULi_4_mult_15_n69) );
  OAI22X1 U826 ( .A0(n487), .A1(n446), .B0(n488), .B1(n447), .Y(
        MULi_4_mult_15_n68) );
  OAI22X1 U827 ( .A0(n485), .A1(n436), .B0(n440), .B1(n486), .Y(
        MULi_4_mult_15_n61) );
  OAI22X1 U828 ( .A0(n487), .A1(n445), .B0(n488), .B1(n446), .Y(
        MULi_4_mult_15_n67) );
  OAI22X1 U829 ( .A0(n485), .A1(n435), .B0(n486), .B1(n436), .Y(
        MULi_4_mult_15_n60) );
  OAI22X1 U830 ( .A0(n487), .A1(n444), .B0(n488), .B1(n445), .Y(
        MULi_4_mult_15_n66) );
  OAI22X1 U831 ( .A0(n487), .A1(n443), .B0(n488), .B1(n444), .Y(
        MULi_4_mult_15_n65) );
  OAI22X1 U832 ( .A0(n485), .A1(n434), .B0(n486), .B1(n435), .Y(
        MULi_4_mult_15_n59) );
  INVX4 U833 ( .A(n78), .Y(n455) );
  AOI22X2 U834 ( .A0(TEMP_H[28]), .A1(n501), .B0(n545), .B1(n534), .Y(n498) );
  AOI22X2 U835 ( .A0(n546), .A1(n539), .B0(TEMP_H[25]), .B1(n512), .Y(n515) );
  AOI22X1 U836 ( .A0(n548), .A1(n538), .B0(TEMP_H[26]), .B1(n152), .Y(n540) );
  AOI22X2 U837 ( .A0(n548), .A1(n539), .B0(TEMP_H[25]), .B1(n152), .Y(n541) );
  AOI22X2 U838 ( .A0(n547), .A1(TEMP_H[31]), .B0(n528), .B1(n524), .Y(n517) );
  OAI21X1 U839 ( .A0(n519), .A1(n171), .B0(n517), .Y(MULi_3_mult_15_n72) );
  AOI22X2 U840 ( .A0(TEMP_H[25]), .A1(n501), .B0(n545), .B1(n539), .Y(n504) );
  AOI22X2 U841 ( .A0(TEMP_H[26]), .A1(n501), .B0(n545), .B1(n538), .Y(n500) );
  AOI22X2 U842 ( .A0(TEMP_H[27]), .A1(n501), .B0(n545), .B1(n536), .Y(n499) );
  OAI22X1 U843 ( .A0(n549), .A1(n496), .B0(n550), .B1(n497), .Y(
        MULi_3_mult_15_n57) );
  OAI22X1 U844 ( .A0(n549), .A1(n497), .B0(n550), .B1(n498), .Y(
        MULi_3_mult_15_n58) );
  OAI22X1 U845 ( .A0(n551), .A1(n515), .B0(n552), .B1(n513), .Y(
        MULi_3_mult_15_n70) );
  OAI22X1 U846 ( .A0(n544), .A1(n540), .B0(n542), .B1(n541), .Y(
        MULi_3_mult_15_n86) );
  AOI21X1 U847 ( .A0(SR_to_MUL[24]), .A1(TEMP_H[24]), .B0(n152), .Y(
        MULi_3_mult_15_n55) );
  OAI22X1 U848 ( .A0(TEMP_H[24]), .A1(n542), .B0(n544), .B1(n541), .Y(
        MULi_3_mult_15_n87) );
  ADDFX1 U849 ( .A(MULi_3_mult_15_n19), .B(MULi_3_mult_15_n18), .CI(
        MULi_3_mult_15_n4), .CO(MULi_3_mult_15_n3), .S(MUL_to_PIPE1[60]) );
  ADDFX1 U850 ( .A(MULi_3_mult_15_n17), .B(MULi_3_mult_15_n16), .CI(
        MULi_3_mult_15_n3), .CO(MULi_3_mult_15_n2), .S(MUL_to_PIPE1[61]) );
  ADDFX1 U851 ( .A(MULi_3_mult_15_n15), .B(MULi_3_mult_15_n56), .CI(
        MULi_3_mult_15_n2), .CO(MULi_3_mult_15_n1), .S(MUL_to_PIPE1[62]) );
  OAI22X1 U852 ( .A0(n549), .A1(n504), .B0(n550), .B1(n502), .Y(
        MULi_3_mult_15_n62) );
  OAI22X1 U853 ( .A0(n551), .A1(n511), .B0(n552), .B1(n515), .Y(
        MULi_3_mult_15_n69) );
  OAI22X1 U854 ( .A0(n551), .A1(n510), .B0(n552), .B1(n511), .Y(
        MULi_3_mult_15_n68) );
  OAI22X1 U855 ( .A0(n549), .A1(n500), .B0(n504), .B1(n550), .Y(
        MULi_3_mult_15_n61) );
  OAI22X1 U856 ( .A0(n551), .A1(n509), .B0(n552), .B1(n510), .Y(
        MULi_3_mult_15_n67) );
  OAI22X1 U857 ( .A0(n549), .A1(n499), .B0(n550), .B1(n500), .Y(
        MULi_3_mult_15_n60) );
  OAI22X1 U858 ( .A0(n551), .A1(n508), .B0(n552), .B1(n509), .Y(
        MULi_3_mult_15_n66) );
  OAI22X1 U859 ( .A0(n551), .A1(n507), .B0(n552), .B1(n508), .Y(
        MULi_3_mult_15_n65) );
  OAI22X1 U860 ( .A0(n549), .A1(n498), .B0(n550), .B1(n499), .Y(
        MULi_3_mult_15_n59) );
  INVX4 U861 ( .A(n74), .Y(n519) );
  AOI22X2 U862 ( .A0(TEMP_H[36]), .A1(n565), .B0(n609), .B1(n598), .Y(n562) );
  AOI22X2 U863 ( .A0(n610), .A1(n603), .B0(TEMP_H[33]), .B1(n576), .Y(n579) );
  AOI22X1 U864 ( .A0(n612), .A1(n602), .B0(TEMP_H[34]), .B1(n153), .Y(n604) );
  AOI22X2 U865 ( .A0(n612), .A1(n603), .B0(TEMP_H[33]), .B1(n153), .Y(n605) );
  AOI22X2 U866 ( .A0(n611), .A1(TEMP_H[39]), .B0(n592), .B1(n588), .Y(n581) );
  OAI21X1 U867 ( .A0(n583), .A1(n173), .B0(n581), .Y(MULi_2_mult_15_n72) );
  AOI22X2 U868 ( .A0(TEMP_H[33]), .A1(n565), .B0(n609), .B1(n603), .Y(n568) );
  AOI22X2 U869 ( .A0(TEMP_H[34]), .A1(n565), .B0(n609), .B1(n602), .Y(n564) );
  AOI22X2 U870 ( .A0(TEMP_H[35]), .A1(n565), .B0(n609), .B1(n600), .Y(n563) );
  OAI22X1 U871 ( .A0(n613), .A1(n560), .B0(n614), .B1(n561), .Y(
        MULi_2_mult_15_n57) );
  OAI22X1 U872 ( .A0(n613), .A1(n561), .B0(n614), .B1(n562), .Y(
        MULi_2_mult_15_n58) );
  OAI22X1 U873 ( .A0(n615), .A1(n579), .B0(n616), .B1(n577), .Y(
        MULi_2_mult_15_n70) );
  OAI22X1 U874 ( .A0(n608), .A1(n604), .B0(n606), .B1(n605), .Y(
        MULi_2_mult_15_n86) );
  AOI21X1 U875 ( .A0(SR_to_MUL[32]), .A1(TEMP_H[32]), .B0(n153), .Y(
        MULi_2_mult_15_n55) );
  OAI22X1 U876 ( .A0(TEMP_H[32]), .A1(n606), .B0(n608), .B1(n605), .Y(
        MULi_2_mult_15_n87) );
  OAI22X1 U877 ( .A0(n613), .A1(n568), .B0(n614), .B1(n566), .Y(
        MULi_2_mult_15_n62) );
  OAI22X1 U878 ( .A0(n615), .A1(n575), .B0(n616), .B1(n579), .Y(
        MULi_2_mult_15_n69) );
  OAI22X1 U879 ( .A0(n615), .A1(n574), .B0(n616), .B1(n575), .Y(
        MULi_2_mult_15_n68) );
  OAI22X1 U880 ( .A0(n613), .A1(n564), .B0(n568), .B1(n614), .Y(
        MULi_2_mult_15_n61) );
  OAI22X1 U881 ( .A0(n615), .A1(n573), .B0(n616), .B1(n574), .Y(
        MULi_2_mult_15_n67) );
  OAI22X1 U882 ( .A0(n613), .A1(n563), .B0(n614), .B1(n564), .Y(
        MULi_2_mult_15_n60) );
  OAI22X1 U883 ( .A0(n615), .A1(n572), .B0(n616), .B1(n573), .Y(
        MULi_2_mult_15_n66) );
  OAI22X1 U884 ( .A0(n615), .A1(n571), .B0(n616), .B1(n572), .Y(
        MULi_2_mult_15_n65) );
  OAI22X1 U885 ( .A0(n613), .A1(n562), .B0(n614), .B1(n563), .Y(
        MULi_2_mult_15_n59) );
  INVX4 U886 ( .A(n77), .Y(n583) );
  AOI22X2 U887 ( .A0(TEMP_H[44]), .A1(n629), .B0(n673), .B1(n662), .Y(n626) );
  AOI22X2 U888 ( .A0(n674), .A1(n667), .B0(TEMP_H[41]), .B1(n640), .Y(n643) );
  AOI22X1 U889 ( .A0(n676), .A1(n666), .B0(TEMP_H[42]), .B1(n148), .Y(n668) );
  AOI22X2 U890 ( .A0(n676), .A1(n667), .B0(TEMP_H[41]), .B1(n148), .Y(n669) );
  AOI22X2 U891 ( .A0(n675), .A1(TEMP_H[47]), .B0(n656), .B1(n652), .Y(n645) );
  OAI21X1 U892 ( .A0(n647), .A1(n175), .B0(n645), .Y(MULi_1_mult_15_n72) );
  AOI22X2 U893 ( .A0(TEMP_H[41]), .A1(n629), .B0(n673), .B1(n667), .Y(n632) );
  AOI22X2 U894 ( .A0(TEMP_H[42]), .A1(n629), .B0(n673), .B1(n666), .Y(n628) );
  AOI22X2 U895 ( .A0(TEMP_H[43]), .A1(n629), .B0(n673), .B1(n664), .Y(n627) );
  OAI22X1 U896 ( .A0(n677), .A1(n624), .B0(n678), .B1(n625), .Y(
        MULi_1_mult_15_n57) );
  OAI22X1 U897 ( .A0(n677), .A1(n625), .B0(n678), .B1(n626), .Y(
        MULi_1_mult_15_n58) );
  OAI22X1 U898 ( .A0(n679), .A1(n643), .B0(n680), .B1(n641), .Y(
        MULi_1_mult_15_n70) );
  OAI22X1 U899 ( .A0(n672), .A1(n668), .B0(n670), .B1(n669), .Y(
        MULi_1_mult_15_n86) );
  AOI21X1 U900 ( .A0(SR_to_MUL[40]), .A1(TEMP_H[40]), .B0(n148), .Y(
        MULi_1_mult_15_n55) );
  OAI22X1 U901 ( .A0(TEMP_H[40]), .A1(n670), .B0(n672), .B1(n669), .Y(
        MULi_1_mult_15_n87) );
  ADDFX1 U902 ( .A(MULi_1_mult_15_n19), .B(MULi_1_mult_15_n18), .CI(
        MULi_1_mult_15_n4), .CO(MULi_1_mult_15_n3), .S(MUL_to_PIPE1[92]) );
  ADDFX1 U903 ( .A(MULi_1_mult_15_n17), .B(MULi_1_mult_15_n16), .CI(
        MULi_1_mult_15_n3), .CO(MULi_1_mult_15_n2), .S(MUL_to_PIPE1[93]) );
  ADDFX1 U904 ( .A(MULi_1_mult_15_n15), .B(MULi_1_mult_15_n56), .CI(
        MULi_1_mult_15_n2), .CO(MULi_1_mult_15_n1), .S(MUL_to_PIPE1[94]) );
  OAI22X1 U905 ( .A0(n677), .A1(n632), .B0(n678), .B1(n630), .Y(
        MULi_1_mult_15_n62) );
  OAI22X1 U906 ( .A0(n679), .A1(n639), .B0(n680), .B1(n643), .Y(
        MULi_1_mult_15_n69) );
  OAI22X1 U907 ( .A0(n679), .A1(n638), .B0(n680), .B1(n639), .Y(
        MULi_1_mult_15_n68) );
  OAI22X1 U908 ( .A0(n677), .A1(n628), .B0(n632), .B1(n678), .Y(
        MULi_1_mult_15_n61) );
  OAI22X1 U909 ( .A0(n679), .A1(n637), .B0(n680), .B1(n638), .Y(
        MULi_1_mult_15_n67) );
  OAI22X1 U910 ( .A0(n677), .A1(n627), .B0(n678), .B1(n628), .Y(
        MULi_1_mult_15_n60) );
  OAI22X1 U911 ( .A0(n679), .A1(n636), .B0(n680), .B1(n637), .Y(
        MULi_1_mult_15_n66) );
  OAI22X1 U912 ( .A0(n679), .A1(n635), .B0(n680), .B1(n636), .Y(
        MULi_1_mult_15_n65) );
  OAI22X1 U913 ( .A0(n677), .A1(n626), .B0(n678), .B1(n627), .Y(
        MULi_1_mult_15_n59) );
  INVX4 U914 ( .A(n75), .Y(n647) );
  OAI2BB1X2 U915 ( .A0N(ADD_esteso_12__1_), .A1N(ADD_esteso_13__1_), .B0(n681), 
        .Y(n682) );
endmodule

