package imem_mau is
   -- created by generatebits
   constant IMEMMAUWIDTH : positive := 42;
end imem_mau;
