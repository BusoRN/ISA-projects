package toplevel_params is
  constant fu_LSU_dataw : integer := 32;
  constant fu_LSU_addrw : integer := 15;
end toplevel_params;
