package testbench_constants is
-- width of the data memory
constant DMEMDATAWIDTH : positive := 32;
-- address width of the data memory
constant DMEMADDRWIDTH : positive := 15-2;
-- simulation run time
constant RUNTIME : time := 10000 ns;
-- memory init files
constant DMEM_INIT_FILE : string := "tb/dmem_init.img";
constant IMEM_INIT_FILE : string := "tb/imem_init.img";
end testbench_constants;
