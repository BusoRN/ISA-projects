
module toplevel ( clk, rstx, busy, imem_en_x, imem_addr, imem_data, pc_init, 
        fu_LSU_data_in, fu_LSU_data_out, fu_LSU_addr, fu_LSU_mem_en_x, 
        fu_LSU_wr_en_x, fu_LSU_wr_mask_x );
  output [14:0] imem_addr;
  input [41:0] imem_data;
  input [14:0] pc_init;
  input [31:0] fu_LSU_data_in;
  output [31:0] fu_LSU_data_out;
  output [12:0] fu_LSU_addr;
  output [0:0] fu_LSU_mem_en_x;
  output [0:0] fu_LSU_wr_en_x;
  output [31:0] fu_LSU_wr_mask_x;
  input clk, rstx, busy;
  output imem_en_x;
  wire   inst_fetch_pc_load_wire, inst_fetch_ra_load_wire,
         inst_fetch_pc_opcode_wire_0_, ic_simm_cntrl_B1_wire_0_,
         ic_socket_lsu_o1_bus_cntrl_wire_0_, ic_socket_RF_o1_bus_cntrl_wire_0_,
         ic_socket_bool_o1_bus_cntrl_wire_0_,
         ic_socket_gcu_o1_bus_cntrl_wire_0_,
         ic_socket_ALU_o1_bus_cntrl_wire_0_,
         ic_socket_LIFTING_o1_bus_cntrl_wire_0_, fu_LSU_t1load_wire,
         fu_LSU_o1load_wire, fu_ALU_t1load_wire, fu_LIFTING_in1_load_wire,
         fu_LIFTING_in2_load_wire, rf_RF_t1load_wire, rf_BOOL_t1load_wire,
         rf_BOOL_t1opcode_wire_0_, rf_BOOL_r1opcode_wire_0_,
         inst_fetch_increased_pc_0_, inst_fetch_increased_pc_1_,
         inst_fetch_increased_pc_2_, inst_fetch_increased_pc_3_,
         inst_fetch_increased_pc_4_, inst_fetch_increased_pc_5_,
         inst_fetch_increased_pc_6_, inst_fetch_increased_pc_7_,
         inst_fetch_increased_pc_8_, inst_fetch_increased_pc_9_,
         inst_fetch_increased_pc_10_, inst_fetch_increased_pc_11_,
         inst_fetch_increased_pc_12_, inst_fetch_increased_pc_13_,
         inst_fetch_increased_pc_14_, inst_fetch_N79, inst_fetch_N76,
         inst_fetch_N75, inst_fetch_N74, inst_fetch_N73, inst_fetch_N72,
         inst_fetch_N71, inst_fetch_N70, inst_fetch_N69, inst_fetch_N68,
         inst_fetch_N67, inst_fetch_N66, inst_fetch_N65, inst_fetch_N64,
         inst_fetch_N63, inst_fetch_N62, inst_fetch_N61, inst_fetch_N60,
         inst_fetch_N59, inst_fetch_N58, inst_fetch_N57, inst_fetch_N56,
         inst_fetch_N55, inst_fetch_N54, inst_fetch_N53, inst_fetch_N52,
         inst_fetch_N51, inst_fetch_N50, inst_fetch_N49, inst_fetch_N48,
         inst_fetch_N47, inst_fetch_reset_cntr_0_, inst_fetch_reset_cntr_1_,
         inst_fetch_reset_cntr_2_, inst_fetch_reset_cntr_3_,
         inst_fetch_reset_cntr_4_, inst_fetch_reset_cntr_5_,
         inst_fetch_reset_cntr_6_, inst_fetch_reset_cntr_7_,
         inst_fetch_reset_cntr_8_, inst_fetch_reset_cntr_9_,
         inst_fetch_reset_cntr_10_, inst_fetch_reset_cntr_11_,
         inst_fetch_reset_cntr_12_, inst_fetch_reset_cntr_13_,
         inst_fetch_reset_cntr_14_, inst_fetch_reset_cntr_15_,
         inst_fetch_reset_cntr_16_, inst_fetch_reset_cntr_17_,
         inst_fetch_reset_cntr_18_, inst_fetch_reset_cntr_19_,
         inst_fetch_reset_cntr_20_, inst_fetch_reset_cntr_21_,
         inst_fetch_reset_cntr_22_, inst_fetch_reset_cntr_23_,
         inst_fetch_reset_cntr_24_, inst_fetch_reset_cntr_25_,
         inst_fetch_reset_cntr_26_, inst_fetch_reset_cntr_27_,
         inst_fetch_reset_cntr_28_, inst_fetch_reset_cntr_29_,
         inst_fetch_reset_cntr_30_, inst_fetch_reset_cntr_31_,
         inst_fetch_reset_lock, inst_fetch_pc_reg_0_, inst_fetch_pc_reg_1_,
         inst_fetch_pc_reg_2_, inst_fetch_pc_reg_3_, inst_fetch_pc_reg_4_,
         inst_fetch_pc_reg_5_, inst_fetch_pc_reg_6_, inst_fetch_pc_reg_7_,
         inst_fetch_pc_reg_8_, inst_fetch_pc_reg_9_, inst_fetch_pc_reg_10_,
         inst_fetch_pc_reg_11_, inst_fetch_pc_reg_12_, inst_fetch_pc_reg_13_,
         inst_fetch_pc_reg_14_, inst_decoder_N232, inst_decoder_N230,
         inst_decoder_N121, inst_decoder_N119, fu_LSU_o1shadow_reg_0_,
         fu_LSU_o1shadow_reg_1_, fu_LSU_o1shadow_reg_2_,
         fu_LSU_o1shadow_reg_3_, fu_LSU_o1shadow_reg_4_,
         fu_LSU_o1shadow_reg_5_, fu_LSU_o1shadow_reg_6_,
         fu_LSU_o1shadow_reg_7_, fu_LSU_o1shadow_reg_8_,
         fu_LSU_o1shadow_reg_9_, fu_LSU_o1shadow_reg_10_,
         fu_LSU_o1shadow_reg_11_, fu_LSU_o1shadow_reg_12_,
         fu_LSU_o1shadow_reg_13_, fu_LSU_o1shadow_reg_14_,
         fu_LSU_o1shadow_reg_15_, fu_LSU_o1shadow_reg_16_,
         fu_LSU_o1shadow_reg_17_, fu_LSU_o1shadow_reg_18_,
         fu_LSU_o1shadow_reg_19_, fu_LSU_o1shadow_reg_20_,
         fu_LSU_o1shadow_reg_21_, fu_LSU_o1shadow_reg_22_,
         fu_LSU_o1shadow_reg_23_, fu_LSU_o1shadow_reg_24_,
         fu_LSU_o1shadow_reg_25_, fu_LSU_o1shadow_reg_26_,
         fu_LSU_o1shadow_reg_27_, fu_LSU_o1shadow_reg_28_,
         fu_LSU_o1shadow_reg_29_, fu_LSU_o1shadow_reg_30_,
         fu_LSU_o1shadow_reg_31_, fu_LSU_status_addr_reg_0__2_,
         fu_LSU_status_addr_reg_1__0_, fu_LSU_status_addr_reg_1__1_,
         fu_LSU_status_addr_reg_1__2_, fu_LSU_status_addr_reg_1__3_,
         fu_LSU_status_addr_reg_1__4_, rf_RF_reg_0__0_, rf_RF_reg_0__1_,
         rf_RF_reg_0__2_, rf_RF_reg_0__3_, rf_RF_reg_0__4_, rf_RF_reg_0__5_,
         rf_RF_reg_0__6_, rf_RF_reg_0__7_, rf_RF_reg_0__8_, rf_RF_reg_0__9_,
         rf_RF_reg_0__10_, rf_RF_reg_0__11_, rf_RF_reg_0__12_,
         rf_RF_reg_0__13_, rf_RF_reg_0__14_, rf_RF_reg_0__15_,
         rf_RF_reg_0__16_, rf_RF_reg_0__17_, rf_RF_reg_0__18_,
         rf_RF_reg_0__19_, rf_RF_reg_0__20_, rf_RF_reg_0__21_,
         rf_RF_reg_0__22_, rf_RF_reg_0__23_, rf_RF_reg_0__24_,
         rf_RF_reg_0__25_, rf_RF_reg_0__26_, rf_RF_reg_0__27_,
         rf_RF_reg_0__28_, rf_RF_reg_0__29_, rf_RF_reg_0__30_,
         rf_RF_reg_0__31_, rf_RF_reg_1__0_, rf_RF_reg_1__1_, rf_RF_reg_1__2_,
         rf_RF_reg_1__3_, rf_RF_reg_1__4_, rf_RF_reg_1__5_, rf_RF_reg_1__6_,
         rf_RF_reg_1__7_, rf_RF_reg_1__8_, rf_RF_reg_1__9_, rf_RF_reg_1__10_,
         rf_RF_reg_1__11_, rf_RF_reg_1__12_, rf_RF_reg_1__13_,
         rf_RF_reg_1__14_, rf_RF_reg_1__15_, rf_RF_reg_1__16_,
         rf_RF_reg_1__17_, rf_RF_reg_1__18_, rf_RF_reg_1__19_,
         rf_RF_reg_1__20_, rf_RF_reg_1__21_, rf_RF_reg_1__22_,
         rf_RF_reg_1__23_, rf_RF_reg_1__24_, rf_RF_reg_1__25_,
         rf_RF_reg_1__26_, rf_RF_reg_1__27_, rf_RF_reg_1__28_,
         rf_RF_reg_1__29_, rf_RF_reg_1__30_, rf_RF_reg_1__31_, rf_RF_reg_2__0_,
         rf_RF_reg_2__1_, rf_RF_reg_2__2_, rf_RF_reg_2__3_, rf_RF_reg_2__4_,
         rf_RF_reg_2__5_, rf_RF_reg_2__6_, rf_RF_reg_2__7_, rf_RF_reg_2__8_,
         rf_RF_reg_2__9_, rf_RF_reg_2__10_, rf_RF_reg_2__11_, rf_RF_reg_2__12_,
         rf_RF_reg_2__13_, rf_RF_reg_2__14_, rf_RF_reg_2__15_,
         rf_RF_reg_2__16_, rf_RF_reg_2__17_, rf_RF_reg_2__18_,
         rf_RF_reg_2__19_, rf_RF_reg_2__20_, rf_RF_reg_2__21_,
         rf_RF_reg_2__22_, rf_RF_reg_2__23_, rf_RF_reg_2__24_,
         rf_RF_reg_2__25_, rf_RF_reg_2__26_, rf_RF_reg_2__27_,
         rf_RF_reg_2__28_, rf_RF_reg_2__29_, rf_RF_reg_2__30_,
         rf_RF_reg_2__31_, rf_RF_reg_3__0_, rf_RF_reg_3__1_, rf_RF_reg_3__2_,
         rf_RF_reg_3__3_, rf_RF_reg_3__4_, rf_RF_reg_3__5_, rf_RF_reg_3__6_,
         rf_RF_reg_3__7_, rf_RF_reg_3__8_, rf_RF_reg_3__9_, rf_RF_reg_3__10_,
         rf_RF_reg_3__11_, rf_RF_reg_3__12_, rf_RF_reg_3__13_,
         rf_RF_reg_3__14_, rf_RF_reg_3__15_, rf_RF_reg_3__16_,
         rf_RF_reg_3__17_, rf_RF_reg_3__18_, rf_RF_reg_3__19_,
         rf_RF_reg_3__20_, rf_RF_reg_3__21_, rf_RF_reg_3__22_,
         rf_RF_reg_3__23_, rf_RF_reg_3__24_, rf_RF_reg_3__25_,
         rf_RF_reg_3__26_, rf_RF_reg_3__27_, rf_RF_reg_3__28_,
         rf_RF_reg_3__29_, rf_RF_reg_3__30_, rf_RF_reg_3__31_, rf_RF_reg_4__0_,
         rf_RF_reg_4__1_, rf_RF_reg_4__2_, rf_RF_reg_4__3_, rf_RF_reg_4__4_,
         rf_RF_reg_4__5_, rf_RF_reg_4__6_, rf_RF_reg_4__7_, rf_RF_reg_4__8_,
         rf_RF_reg_4__9_, rf_RF_reg_4__10_, rf_RF_reg_4__11_, rf_RF_reg_4__12_,
         rf_RF_reg_4__13_, rf_RF_reg_4__14_, rf_RF_reg_4__15_,
         rf_RF_reg_4__16_, rf_RF_reg_4__17_, rf_RF_reg_4__18_,
         rf_RF_reg_4__19_, rf_RF_reg_4__20_, rf_RF_reg_4__21_,
         rf_RF_reg_4__22_, rf_RF_reg_4__23_, rf_RF_reg_4__24_,
         rf_RF_reg_4__25_, rf_RF_reg_4__26_, rf_RF_reg_4__27_,
         rf_RF_reg_4__28_, rf_RF_reg_4__29_, rf_RF_reg_4__30_,
         rf_RF_reg_4__31_, rf_BOOL_reg_0__0_, rf_BOOL_reg_1__0_, n19, n20, n21,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n43, n44, n45, n46, n47, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n239, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n272, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n408, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n426, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n588, n589, n590, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n625,
         n626, n627, n628, n629, n630, n631, n632, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, fu_ALU_fu_arch_n767, fu_ALU_fu_arch_n766,
         fu_ALU_fu_arch_n765, fu_ALU_fu_arch_n764, fu_ALU_fu_arch_n763,
         fu_ALU_fu_arch_n762, fu_ALU_fu_arch_n761, fu_ALU_fu_arch_n760,
         fu_ALU_fu_arch_n759, fu_ALU_fu_arch_n758, fu_ALU_fu_arch_n757,
         fu_ALU_fu_arch_n756, fu_ALU_fu_arch_n755, fu_ALU_fu_arch_n754,
         fu_ALU_fu_arch_n753, fu_ALU_fu_arch_n752, fu_ALU_fu_arch_n751,
         fu_ALU_fu_arch_n750, fu_ALU_fu_arch_n748, fu_ALU_fu_arch_n747,
         fu_ALU_fu_arch_n746, fu_ALU_fu_arch_n745, fu_ALU_fu_arch_n744,
         fu_ALU_fu_arch_n743, fu_ALU_fu_arch_n742, fu_ALU_fu_arch_n741,
         fu_ALU_fu_arch_n740, fu_ALU_fu_arch_n739, fu_ALU_fu_arch_n738,
         fu_ALU_fu_arch_n737, fu_ALU_fu_arch_n736, fu_ALU_fu_arch_n735,
         fu_ALU_fu_arch_n734, fu_ALU_fu_arch_n733, fu_ALU_fu_arch_n732,
         fu_ALU_fu_arch_n731, fu_ALU_fu_arch_n730, fu_ALU_fu_arch_n729,
         fu_ALU_fu_arch_n728, fu_ALU_fu_arch_n727, fu_ALU_fu_arch_n726,
         fu_ALU_fu_arch_n725, fu_ALU_fu_arch_n724, fu_ALU_fu_arch_n723,
         fu_ALU_fu_arch_n722, fu_ALU_fu_arch_n721, fu_ALU_fu_arch_n720,
         fu_ALU_fu_arch_n719, fu_ALU_fu_arch_n718, fu_ALU_fu_arch_n717,
         fu_ALU_fu_arch_n716, fu_ALU_fu_arch_n715, fu_ALU_fu_arch_n714,
         fu_ALU_fu_arch_n713, fu_ALU_fu_arch_n712, fu_ALU_fu_arch_n711,
         fu_ALU_fu_arch_n710, fu_ALU_fu_arch_n709, fu_ALU_fu_arch_n708,
         fu_ALU_fu_arch_n707, fu_ALU_fu_arch_n706, fu_ALU_fu_arch_n705,
         fu_ALU_fu_arch_n704, fu_ALU_fu_arch_n703, fu_ALU_fu_arch_n702,
         fu_ALU_fu_arch_n701, fu_ALU_fu_arch_n699, fu_ALU_fu_arch_n698,
         fu_ALU_fu_arch_n697, fu_ALU_fu_arch_n696, fu_ALU_fu_arch_n695,
         fu_ALU_fu_arch_n694, fu_ALU_fu_arch_n693, fu_ALU_fu_arch_n692,
         fu_ALU_fu_arch_n691, fu_ALU_fu_arch_n690, fu_ALU_fu_arch_n689,
         fu_ALU_fu_arch_n688, fu_ALU_fu_arch_n687, fu_ALU_fu_arch_n686,
         fu_ALU_fu_arch_n685, fu_ALU_fu_arch_n683, fu_ALU_fu_arch_n682,
         fu_ALU_fu_arch_n681, fu_ALU_fu_arch_n680, fu_ALU_fu_arch_n679,
         fu_ALU_fu_arch_n678, fu_ALU_fu_arch_n677, fu_ALU_fu_arch_n676,
         fu_ALU_fu_arch_n675, fu_ALU_fu_arch_n674, fu_ALU_fu_arch_n673,
         fu_ALU_fu_arch_n672, fu_ALU_fu_arch_n671, fu_ALU_fu_arch_n670,
         fu_ALU_fu_arch_n669, fu_ALU_fu_arch_n668, fu_ALU_fu_arch_n667,
         fu_ALU_fu_arch_n666, fu_ALU_fu_arch_n665, fu_ALU_fu_arch_n664,
         fu_ALU_fu_arch_n663, fu_ALU_fu_arch_n662, fu_ALU_fu_arch_n661,
         fu_ALU_fu_arch_n660, fu_ALU_fu_arch_n659, fu_ALU_fu_arch_n658,
         fu_ALU_fu_arch_n657, fu_ALU_fu_arch_n656, fu_ALU_fu_arch_n655,
         fu_ALU_fu_arch_n654, fu_ALU_fu_arch_n653, fu_ALU_fu_arch_n652,
         fu_ALU_fu_arch_n651, fu_ALU_fu_arch_n650, fu_ALU_fu_arch_n649,
         fu_ALU_fu_arch_n648, fu_ALU_fu_arch_n647, fu_ALU_fu_arch_n645,
         fu_ALU_fu_arch_n644, fu_ALU_fu_arch_n643, fu_ALU_fu_arch_n642,
         fu_ALU_fu_arch_n641, fu_ALU_fu_arch_n640, fu_ALU_fu_arch_n639,
         fu_ALU_fu_arch_n638, fu_ALU_fu_arch_n637, fu_ALU_fu_arch_n636,
         fu_ALU_fu_arch_n635, fu_ALU_fu_arch_n634, fu_ALU_fu_arch_n633,
         fu_ALU_fu_arch_n631, fu_ALU_fu_arch_n630, fu_ALU_fu_arch_n629,
         fu_ALU_fu_arch_n628, fu_ALU_fu_arch_n627, fu_ALU_fu_arch_n626,
         fu_ALU_fu_arch_n625, fu_ALU_fu_arch_n624, fu_ALU_fu_arch_n623,
         fu_ALU_fu_arch_n622, fu_ALU_fu_arch_n621, fu_ALU_fu_arch_n620,
         fu_ALU_fu_arch_n619, fu_ALU_fu_arch_n618, fu_ALU_fu_arch_n617,
         fu_ALU_fu_arch_n616, fu_ALU_fu_arch_n615, fu_ALU_fu_arch_n614,
         fu_ALU_fu_arch_n613, fu_ALU_fu_arch_n612, fu_ALU_fu_arch_n611,
         fu_ALU_fu_arch_n610, fu_ALU_fu_arch_n609, fu_ALU_fu_arch_n608,
         fu_ALU_fu_arch_n607, fu_ALU_fu_arch_n606, fu_ALU_fu_arch_n605,
         fu_ALU_fu_arch_n604, fu_ALU_fu_arch_n603, fu_ALU_fu_arch_n602,
         fu_ALU_fu_arch_n601, fu_ALU_fu_arch_n600, fu_ALU_fu_arch_n599,
         fu_ALU_fu_arch_n598, fu_ALU_fu_arch_n596, fu_ALU_fu_arch_n595,
         fu_ALU_fu_arch_n594, fu_ALU_fu_arch_n593, fu_ALU_fu_arch_n592,
         fu_ALU_fu_arch_n591, fu_ALU_fu_arch_n590, fu_ALU_fu_arch_n589,
         fu_ALU_fu_arch_n588, fu_ALU_fu_arch_n587, fu_ALU_fu_arch_n586,
         fu_ALU_fu_arch_n585, fu_ALU_fu_arch_n584, fu_ALU_fu_arch_n583,
         fu_ALU_fu_arch_n581, fu_ALU_fu_arch_n580, fu_ALU_fu_arch_n579,
         fu_ALU_fu_arch_n578, fu_ALU_fu_arch_n577, fu_ALU_fu_arch_n575,
         fu_ALU_fu_arch_n574, fu_ALU_fu_arch_n573, fu_ALU_fu_arch_n572,
         fu_ALU_fu_arch_n571, fu_ALU_fu_arch_n570, fu_ALU_fu_arch_n569,
         fu_ALU_fu_arch_n568, fu_ALU_fu_arch_n567, fu_ALU_fu_arch_n566,
         fu_ALU_fu_arch_n564, fu_ALU_fu_arch_n563, fu_ALU_fu_arch_n562,
         fu_ALU_fu_arch_n561, fu_ALU_fu_arch_n560, fu_ALU_fu_arch_n559,
         fu_ALU_fu_arch_n556, fu_ALU_fu_arch_n555, fu_ALU_fu_arch_n554,
         fu_ALU_fu_arch_n553, fu_ALU_fu_arch_n552, fu_ALU_fu_arch_n551,
         fu_ALU_fu_arch_n550, fu_ALU_fu_arch_n549, fu_ALU_fu_arch_n548,
         fu_ALU_fu_arch_n547, fu_ALU_fu_arch_n546, fu_ALU_fu_arch_n545,
         fu_ALU_fu_arch_n544, fu_ALU_fu_arch_n543, fu_ALU_fu_arch_n542,
         fu_ALU_fu_arch_n541, fu_ALU_fu_arch_n540, fu_ALU_fu_arch_n539,
         fu_ALU_fu_arch_n538, fu_ALU_fu_arch_n537, fu_ALU_fu_arch_n536,
         fu_ALU_fu_arch_n535, fu_ALU_fu_arch_n534, fu_ALU_fu_arch_n533,
         fu_ALU_fu_arch_n532, fu_ALU_fu_arch_n531, fu_ALU_fu_arch_n530,
         fu_ALU_fu_arch_n529, fu_ALU_fu_arch_n528, fu_ALU_fu_arch_n527,
         fu_ALU_fu_arch_n526, fu_ALU_fu_arch_n525, fu_ALU_fu_arch_n524,
         fu_ALU_fu_arch_n523, fu_ALU_fu_arch_n522, fu_ALU_fu_arch_n521,
         fu_ALU_fu_arch_n520, fu_ALU_fu_arch_n519, fu_ALU_fu_arch_n518,
         fu_ALU_fu_arch_n517, fu_ALU_fu_arch_n516, fu_ALU_fu_arch_n515,
         fu_ALU_fu_arch_n514, fu_ALU_fu_arch_n513, fu_ALU_fu_arch_n512,
         fu_ALU_fu_arch_n511, fu_ALU_fu_arch_n510, fu_ALU_fu_arch_n509,
         fu_ALU_fu_arch_n508, fu_ALU_fu_arch_n507, fu_ALU_fu_arch_n506,
         fu_ALU_fu_arch_n505, fu_ALU_fu_arch_n504, fu_ALU_fu_arch_n503,
         fu_ALU_fu_arch_n502, fu_ALU_fu_arch_n501, fu_ALU_fu_arch_n500,
         fu_ALU_fu_arch_n499, fu_ALU_fu_arch_n498, fu_ALU_fu_arch_n497,
         fu_ALU_fu_arch_n496, fu_ALU_fu_arch_n495, fu_ALU_fu_arch_n494,
         fu_ALU_fu_arch_n493, fu_ALU_fu_arch_n492, fu_ALU_fu_arch_n491,
         fu_ALU_fu_arch_n490, fu_ALU_fu_arch_n489, fu_ALU_fu_arch_n488,
         fu_ALU_fu_arch_n487, fu_ALU_fu_arch_n486, fu_ALU_fu_arch_n485,
         fu_ALU_fu_arch_n484, fu_ALU_fu_arch_n483, fu_ALU_fu_arch_n482,
         fu_ALU_fu_arch_n481, fu_ALU_fu_arch_n480, fu_ALU_fu_arch_n479,
         fu_ALU_fu_arch_n478, fu_ALU_fu_arch_n477, fu_ALU_fu_arch_n476,
         fu_ALU_fu_arch_n475, fu_ALU_fu_arch_n474, fu_ALU_fu_arch_n473,
         fu_ALU_fu_arch_n472, fu_ALU_fu_arch_n471, fu_ALU_fu_arch_n470,
         fu_ALU_fu_arch_n469, fu_ALU_fu_arch_n468, fu_ALU_fu_arch_n467,
         fu_ALU_fu_arch_n466, fu_ALU_fu_arch_n465, fu_ALU_fu_arch_n464,
         fu_ALU_fu_arch_n463, fu_ALU_fu_arch_n462, fu_ALU_fu_arch_n461,
         fu_ALU_fu_arch_n460, fu_ALU_fu_arch_n459, fu_ALU_fu_arch_n458,
         fu_ALU_fu_arch_n457, fu_ALU_fu_arch_n456, fu_ALU_fu_arch_n455,
         fu_ALU_fu_arch_n454, fu_ALU_fu_arch_n453, fu_ALU_fu_arch_n452,
         fu_ALU_fu_arch_n451, fu_ALU_fu_arch_n450, fu_ALU_fu_arch_n449,
         fu_ALU_fu_arch_n448, fu_ALU_fu_arch_n447, fu_ALU_fu_arch_n446,
         fu_ALU_fu_arch_n445, fu_ALU_fu_arch_n443, fu_ALU_fu_arch_n442,
         fu_ALU_fu_arch_n441, fu_ALU_fu_arch_n440, fu_ALU_fu_arch_n439,
         fu_ALU_fu_arch_n438, fu_ALU_fu_arch_n437, fu_ALU_fu_arch_n436,
         fu_ALU_fu_arch_n435, fu_ALU_fu_arch_n434, fu_ALU_fu_arch_n433,
         fu_ALU_fu_arch_n432, fu_ALU_fu_arch_n431, fu_ALU_fu_arch_n430,
         fu_ALU_fu_arch_n429, fu_ALU_fu_arch_n428, fu_ALU_fu_arch_n427,
         fu_ALU_fu_arch_n425, fu_ALU_fu_arch_n424, fu_ALU_fu_arch_n423,
         fu_ALU_fu_arch_n422, fu_ALU_fu_arch_n421, fu_ALU_fu_arch_n419,
         fu_ALU_fu_arch_n418, fu_ALU_fu_arch_n417, fu_ALU_fu_arch_n416,
         fu_ALU_fu_arch_n415, fu_ALU_fu_arch_n414, fu_ALU_fu_arch_n413,
         fu_ALU_fu_arch_n412, fu_ALU_fu_arch_n411, fu_ALU_fu_arch_n410,
         fu_ALU_fu_arch_n409, fu_ALU_fu_arch_n408, fu_ALU_fu_arch_n407,
         fu_ALU_fu_arch_n406, fu_ALU_fu_arch_n405, fu_ALU_fu_arch_n404,
         fu_ALU_fu_arch_n403, fu_ALU_fu_arch_n400, fu_ALU_fu_arch_n399,
         fu_ALU_fu_arch_n398, fu_ALU_fu_arch_n397, fu_ALU_fu_arch_n396,
         fu_ALU_fu_arch_n395, fu_ALU_fu_arch_n394, fu_ALU_fu_arch_n393,
         fu_ALU_fu_arch_n392, fu_ALU_fu_arch_n391, fu_ALU_fu_arch_n390,
         fu_ALU_fu_arch_n389, fu_ALU_fu_arch_n388, fu_ALU_fu_arch_n387,
         fu_ALU_fu_arch_n386, fu_ALU_fu_arch_n385, fu_ALU_fu_arch_n384,
         fu_ALU_fu_arch_n383, fu_ALU_fu_arch_n382, fu_ALU_fu_arch_n379,
         fu_ALU_fu_arch_n378, fu_ALU_fu_arch_n376, fu_ALU_fu_arch_n374,
         fu_ALU_fu_arch_n373, fu_ALU_fu_arch_n372, fu_ALU_fu_arch_n371,
         fu_ALU_fu_arch_n370, fu_ALU_fu_arch_n369, fu_ALU_fu_arch_n368,
         fu_ALU_fu_arch_n367, fu_ALU_fu_arch_n366, fu_ALU_fu_arch_n365,
         fu_ALU_fu_arch_n364, fu_ALU_fu_arch_n363, fu_ALU_fu_arch_n362,
         fu_ALU_fu_arch_n361, fu_ALU_fu_arch_n360, fu_ALU_fu_arch_n359,
         fu_ALU_fu_arch_n358, fu_ALU_fu_arch_n356, fu_ALU_fu_arch_n354,
         fu_ALU_fu_arch_n353, fu_ALU_fu_arch_n352, fu_ALU_fu_arch_n351,
         fu_ALU_fu_arch_n350, fu_ALU_fu_arch_n349, fu_ALU_fu_arch_n348,
         fu_ALU_fu_arch_n347, fu_ALU_fu_arch_n346, fu_ALU_fu_arch_n345,
         fu_ALU_fu_arch_n344, fu_ALU_fu_arch_n343, fu_ALU_fu_arch_n342,
         fu_ALU_fu_arch_n341, fu_ALU_fu_arch_n340, fu_ALU_fu_arch_n339,
         fu_ALU_fu_arch_n338, fu_ALU_fu_arch_n337, fu_ALU_fu_arch_n336,
         fu_ALU_fu_arch_n335, fu_ALU_fu_arch_n334, fu_ALU_fu_arch_n333,
         fu_ALU_fu_arch_n332, fu_ALU_fu_arch_n331, fu_ALU_fu_arch_n330,
         fu_ALU_fu_arch_n329, fu_ALU_fu_arch_n328, fu_ALU_fu_arch_n327,
         fu_ALU_fu_arch_n326, fu_ALU_fu_arch_n325, fu_ALU_fu_arch_n323,
         fu_ALU_fu_arch_n322, fu_ALU_fu_arch_n321, fu_ALU_fu_arch_n320,
         fu_ALU_fu_arch_n319, fu_ALU_fu_arch_n318, fu_ALU_fu_arch_n317,
         fu_ALU_fu_arch_n316, fu_ALU_fu_arch_n315, fu_ALU_fu_arch_n314,
         fu_ALU_fu_arch_n313, fu_ALU_fu_arch_n312, fu_ALU_fu_arch_n311,
         fu_ALU_fu_arch_n310, fu_ALU_fu_arch_n309, fu_ALU_fu_arch_n308,
         fu_ALU_fu_arch_n307, fu_ALU_fu_arch_n306, fu_ALU_fu_arch_n305,
         fu_ALU_fu_arch_n304, fu_ALU_fu_arch_n303, fu_ALU_fu_arch_n301,
         fu_ALU_fu_arch_n300, fu_ALU_fu_arch_n299, fu_ALU_fu_arch_n298,
         fu_ALU_fu_arch_n297, fu_ALU_fu_arch_n296, fu_ALU_fu_arch_n295,
         fu_ALU_fu_arch_n294, fu_ALU_fu_arch_n293, fu_ALU_fu_arch_n292,
         fu_ALU_fu_arch_n291, fu_ALU_fu_arch_n290, fu_ALU_fu_arch_n289,
         fu_ALU_fu_arch_n288, fu_ALU_fu_arch_n287, fu_ALU_fu_arch_n285,
         fu_ALU_fu_arch_n284, fu_ALU_fu_arch_n283, fu_ALU_fu_arch_n282,
         fu_ALU_fu_arch_n281, fu_ALU_fu_arch_n279, fu_ALU_fu_arch_n278,
         fu_ALU_fu_arch_n277, fu_ALU_fu_arch_n276, fu_ALU_fu_arch_n275,
         fu_ALU_fu_arch_n274, fu_ALU_fu_arch_n271, fu_ALU_fu_arch_n270,
         fu_ALU_fu_arch_n268, fu_ALU_fu_arch_n267, fu_ALU_fu_arch_n266,
         fu_ALU_fu_arch_n265, fu_ALU_fu_arch_n264, fu_ALU_fu_arch_n263,
         fu_ALU_fu_arch_n262, fu_ALU_fu_arch_n260, fu_ALU_fu_arch_n259,
         fu_ALU_fu_arch_n256, fu_ALU_fu_arch_n255, fu_ALU_fu_arch_n254,
         fu_ALU_fu_arch_n253, fu_ALU_fu_arch_n251, fu_ALU_fu_arch_n250,
         fu_ALU_fu_arch_n249, fu_ALU_fu_arch_n248, fu_ALU_fu_arch_n247,
         fu_ALU_fu_arch_n246, fu_ALU_fu_arch_n245, fu_ALU_fu_arch_n243,
         fu_ALU_fu_arch_n242, fu_ALU_fu_arch_n241, fu_ALU_fu_arch_n240,
         fu_ALU_fu_arch_n239, fu_ALU_fu_arch_n236, fu_ALU_fu_arch_n235,
         fu_ALU_fu_arch_n234, fu_ALU_fu_arch_n233, fu_ALU_fu_arch_n232,
         fu_ALU_fu_arch_n231, fu_ALU_fu_arch_n230, fu_ALU_fu_arch_n229,
         fu_ALU_fu_arch_n228, fu_ALU_fu_arch_n227, fu_ALU_fu_arch_n226,
         fu_ALU_fu_arch_n225, fu_ALU_fu_arch_n224, fu_ALU_fu_arch_n223,
         fu_ALU_fu_arch_n221, fu_ALU_fu_arch_n220, fu_ALU_fu_arch_n219,
         fu_ALU_fu_arch_n218, fu_ALU_fu_arch_n217, fu_ALU_fu_arch_n216,
         fu_ALU_fu_arch_n215, fu_ALU_fu_arch_n214, fu_ALU_fu_arch_n213,
         fu_ALU_fu_arch_n212, fu_ALU_fu_arch_n211, fu_ALU_fu_arch_n210,
         fu_ALU_fu_arch_n209, fu_ALU_fu_arch_n208, fu_ALU_fu_arch_n205,
         fu_ALU_fu_arch_n204, fu_ALU_fu_arch_n203, fu_ALU_fu_arch_n202,
         fu_ALU_fu_arch_n201, fu_ALU_fu_arch_n200, fu_ALU_fu_arch_n199,
         fu_ALU_fu_arch_n197, fu_ALU_fu_arch_n196, fu_ALU_fu_arch_n195,
         fu_ALU_fu_arch_n194, fu_ALU_fu_arch_n193, fu_ALU_fu_arch_n192,
         fu_ALU_fu_arch_n191, fu_ALU_fu_arch_n190, fu_ALU_fu_arch_n189,
         fu_ALU_fu_arch_n187, fu_ALU_fu_arch_n186, fu_ALU_fu_arch_n185,
         fu_ALU_fu_arch_n184, fu_ALU_fu_arch_n183, fu_ALU_fu_arch_n182,
         fu_ALU_fu_arch_n181, fu_ALU_fu_arch_n180, fu_ALU_fu_arch_n179,
         fu_ALU_fu_arch_n178, fu_ALU_fu_arch_n177, fu_ALU_fu_arch_n176,
         fu_ALU_fu_arch_n175, fu_ALU_fu_arch_n172, fu_ALU_fu_arch_n171,
         fu_ALU_fu_arch_n170, fu_ALU_fu_arch_n169, fu_ALU_fu_arch_n168,
         fu_ALU_fu_arch_n167, fu_ALU_fu_arch_n166, fu_ALU_fu_arch_n165,
         fu_ALU_fu_arch_n164, fu_ALU_fu_arch_n162, fu_ALU_fu_arch_n160,
         fu_ALU_fu_arch_n159, fu_ALU_fu_arch_n158, fu_ALU_fu_arch_n157,
         fu_ALU_fu_arch_n156, fu_ALU_fu_arch_n155, fu_ALU_fu_arch_n154,
         fu_ALU_fu_arch_n153, fu_ALU_fu_arch_n152, fu_ALU_fu_arch_n151,
         fu_ALU_fu_arch_n148, fu_ALU_fu_arch_n147, fu_ALU_fu_arch_n146,
         fu_ALU_fu_arch_n145, fu_ALU_fu_arch_n144, fu_ALU_fu_arch_n143,
         fu_ALU_fu_arch_n142, fu_ALU_fu_arch_n141, fu_ALU_fu_arch_n140,
         fu_ALU_fu_arch_n139, fu_ALU_fu_arch_n138, fu_ALU_fu_arch_n137,
         fu_ALU_fu_arch_n136, fu_ALU_fu_arch_n135, fu_ALU_fu_arch_n134,
         fu_ALU_fu_arch_n133, fu_ALU_fu_arch_n132, fu_ALU_fu_arch_n131,
         fu_ALU_fu_arch_n130, fu_ALU_fu_arch_n129, fu_ALU_fu_arch_n128,
         fu_ALU_fu_arch_n127, fu_ALU_fu_arch_n126, fu_ALU_fu_arch_n125,
         fu_ALU_fu_arch_n121, fu_ALU_fu_arch_n119, fu_ALU_fu_arch_n118,
         fu_ALU_fu_arch_n117, fu_ALU_fu_arch_n116, fu_ALU_fu_arch_n115,
         fu_ALU_fu_arch_n114, fu_ALU_fu_arch_n113, fu_ALU_fu_arch_n112,
         fu_ALU_fu_arch_n111, fu_ALU_fu_arch_n110, fu_ALU_fu_arch_n109,
         fu_ALU_fu_arch_n108, fu_ALU_fu_arch_n107, fu_ALU_fu_arch_N643,
         fu_ALU_fu_arch_N642, fu_ALU_fu_arch_N641, fu_ALU_fu_arch_N640,
         fu_ALU_fu_arch_N639, fu_ALU_fu_arch_N638, fu_ALU_fu_arch_N637,
         fu_ALU_fu_arch_N636, fu_ALU_fu_arch_N635, fu_ALU_fu_arch_N634,
         fu_ALU_fu_arch_N633, fu_ALU_fu_arch_N632, fu_ALU_fu_arch_N631,
         fu_ALU_fu_arch_N630, fu_ALU_fu_arch_N629, fu_ALU_fu_arch_N628,
         fu_ALU_fu_arch_N627, fu_ALU_fu_arch_N626, fu_ALU_fu_arch_N625,
         fu_ALU_fu_arch_N624, fu_ALU_fu_arch_N623, fu_ALU_fu_arch_N622,
         fu_ALU_fu_arch_N621, fu_ALU_fu_arch_N620, fu_ALU_fu_arch_N619,
         fu_ALU_fu_arch_N618, fu_ALU_fu_arch_N617, fu_ALU_fu_arch_N616,
         fu_ALU_fu_arch_N615, fu_ALU_fu_arch_N614, fu_ALU_fu_arch_N613,
         fu_ALU_fu_arch_N612, fu_ALU_fu_arch_N99, fu_ALU_fu_arch_N98,
         fu_ALU_fu_arch_N97, fu_ALU_fu_arch_N64, fu_ALU_fu_arch_N63,
         fu_ALU_fu_arch_N62, fu_ALU_fu_arch_N61, fu_ALU_fu_arch_N60,
         fu_ALU_fu_arch_N59, fu_ALU_fu_arch_N58, fu_ALU_fu_arch_N57,
         fu_ALU_fu_arch_N56, fu_ALU_fu_arch_N55, fu_ALU_fu_arch_N54,
         fu_ALU_fu_arch_N53, fu_ALU_fu_arch_N52, fu_ALU_fu_arch_N51,
         fu_ALU_fu_arch_N50, fu_ALU_fu_arch_N49, fu_ALU_fu_arch_N48,
         fu_ALU_fu_arch_N47, fu_ALU_fu_arch_N46, fu_ALU_fu_arch_N45,
         fu_ALU_fu_arch_N44, fu_ALU_fu_arch_N43, fu_ALU_fu_arch_N42,
         fu_ALU_fu_arch_N41, fu_ALU_fu_arch_N40, fu_ALU_fu_arch_N39,
         fu_ALU_fu_arch_N38, fu_ALU_fu_arch_N37, fu_ALU_fu_arch_N36,
         fu_ALU_fu_arch_N35, fu_ALU_fu_arch_N34, fu_ALU_fu_arch_N33,
         inst_fetch_add_136_carry_2_, inst_fetch_add_136_carry_3_,
         inst_fetch_add_136_carry_4_, inst_fetch_add_136_carry_5_,
         inst_fetch_add_136_carry_6_, inst_fetch_add_136_carry_7_,
         inst_fetch_add_136_carry_8_, inst_fetch_add_136_carry_9_,
         inst_fetch_add_136_carry_10_, inst_fetch_add_136_carry_11_,
         inst_fetch_add_136_carry_12_, inst_fetch_add_136_carry_13_,
         inst_fetch_add_136_carry_14_, inst_fetch_add_113_carry_2_,
         inst_fetch_add_113_carry_3_, inst_fetch_add_113_carry_4_,
         inst_fetch_add_113_carry_5_, inst_fetch_add_113_carry_6_,
         inst_fetch_add_113_carry_7_, inst_fetch_add_113_carry_8_,
         inst_fetch_add_113_carry_9_, inst_fetch_add_113_carry_10_,
         inst_fetch_add_113_carry_11_, inst_fetch_add_113_carry_12_,
         inst_fetch_add_113_carry_13_, inst_fetch_add_113_carry_14_,
         inst_fetch_add_113_carry_15_, inst_fetch_add_113_carry_16_,
         inst_fetch_add_113_carry_17_, inst_fetch_add_113_carry_18_,
         inst_fetch_add_113_carry_19_, inst_fetch_add_113_carry_20_,
         inst_fetch_add_113_carry_21_, inst_fetch_add_113_carry_22_,
         inst_fetch_add_113_carry_23_, inst_fetch_add_113_carry_24_,
         inst_fetch_add_113_carry_25_, inst_fetch_add_113_carry_26_,
         inst_fetch_add_113_carry_27_, inst_fetch_add_113_carry_28_,
         inst_fetch_add_113_carry_29_, inst_fetch_add_113_carry_30_,
         inst_fetch_add_113_carry_31_, fu_ALU_fu_arch_sub_200_B_not_0_,
         fu_ALU_fu_arch_sub_200_B_not_2_, fu_ALU_fu_arch_sub_200_B_not_4_,
         fu_ALU_fu_arch_sub_200_B_not_6_, fu_ALU_fu_arch_sub_200_B_not_12_,
         fu_ALU_fu_arch_sub_200_B_not_16_, fu_ALU_fu_arch_sub_200_B_not_17_,
         fu_ALU_fu_arch_sub_200_B_not_20_, fu_ALU_fu_arch_sub_200_B_not_21_,
         fu_ALU_fu_arch_sub_200_B_not_22_, fu_ALU_fu_arch_sub_200_B_not_23_,
         fu_ALU_fu_arch_sub_200_B_not_24_, fu_ALU_fu_arch_sub_200_B_not_30_,
         fu_ALU_fu_arch_sub_200_carry_1_, fu_ALU_fu_arch_sub_200_carry_2_,
         fu_ALU_fu_arch_sub_200_carry_3_, fu_ALU_fu_arch_sub_200_carry_4_,
         fu_ALU_fu_arch_sub_200_carry_5_, fu_ALU_fu_arch_sub_200_carry_6_,
         fu_ALU_fu_arch_sub_200_carry_7_, fu_ALU_fu_arch_sub_200_carry_8_,
         fu_ALU_fu_arch_sub_200_carry_9_, fu_ALU_fu_arch_sub_200_carry_10_,
         fu_ALU_fu_arch_sub_200_carry_11_, fu_ALU_fu_arch_sub_200_carry_12_,
         fu_ALU_fu_arch_sub_200_carry_13_, fu_ALU_fu_arch_sub_200_carry_14_,
         fu_ALU_fu_arch_sub_200_carry_15_, fu_ALU_fu_arch_sub_200_carry_16_,
         fu_ALU_fu_arch_sub_200_carry_17_, fu_ALU_fu_arch_sub_200_carry_18_,
         fu_ALU_fu_arch_sub_200_carry_19_, fu_ALU_fu_arch_sub_200_carry_20_,
         fu_ALU_fu_arch_sub_200_carry_21_, fu_ALU_fu_arch_sub_200_carry_22_,
         fu_ALU_fu_arch_sub_200_carry_23_, fu_ALU_fu_arch_sub_200_carry_24_,
         fu_ALU_fu_arch_sub_200_carry_25_, fu_ALU_fu_arch_sub_200_carry_26_,
         fu_ALU_fu_arch_sub_200_carry_27_, fu_ALU_fu_arch_sub_200_carry_28_,
         fu_ALU_fu_arch_sub_200_carry_29_, fu_ALU_fu_arch_sub_200_carry_30_,
         fu_ALU_fu_arch_sub_200_carry_31_, fu_ALU_fu_arch_sub_200_B_2_,
         fu_ALU_fu_arch_sub_200_B_4_, fu_ALU_fu_arch_sub_200_B_5_,
         fu_ALU_fu_arch_sub_200_B_8_, fu_ALU_fu_arch_sub_200_B_9_,
         fu_ALU_fu_arch_sub_200_B_11_, fu_ALU_fu_arch_sub_200_B_14_,
         fu_ALU_fu_arch_sub_200_B_18_, fu_ALU_fu_arch_sub_200_B_19_,
         fu_ALU_fu_arch_sub_200_B_21_, fu_ALU_fu_arch_sub_200_B_22_,
         fu_ALU_fu_arch_sub_200_B_27_, fu_ALU_fu_arch_sub_200_B_29_,
         fu_ALU_fu_arch_sub_200_B_30_, fu_ALU_fu_arch_sub_200_A_1_,
         fu_ALU_fu_arch_lt_gt_188_A_28_, fu_ALU_fu_arch_add_171_carry_1_,
         fu_ALU_fu_arch_add_171_carry_2_, fu_ALU_fu_arch_add_171_carry_3_,
         fu_ALU_fu_arch_add_171_carry_4_, fu_ALU_fu_arch_add_171_carry_5_,
         fu_ALU_fu_arch_add_171_carry_6_, fu_ALU_fu_arch_add_171_carry_7_,
         fu_ALU_fu_arch_add_171_carry_8_, fu_ALU_fu_arch_add_171_carry_9_,
         fu_ALU_fu_arch_add_171_carry_10_, fu_ALU_fu_arch_add_171_carry_11_,
         fu_ALU_fu_arch_add_171_carry_12_, fu_ALU_fu_arch_add_171_carry_13_,
         fu_ALU_fu_arch_add_171_carry_14_, fu_ALU_fu_arch_add_171_carry_15_,
         fu_ALU_fu_arch_add_171_carry_16_, fu_ALU_fu_arch_add_171_carry_17_,
         fu_ALU_fu_arch_add_171_carry_18_, fu_ALU_fu_arch_add_171_carry_19_,
         fu_ALU_fu_arch_add_171_carry_20_, fu_ALU_fu_arch_add_171_carry_21_,
         fu_ALU_fu_arch_add_171_carry_22_, fu_ALU_fu_arch_add_171_carry_23_,
         fu_ALU_fu_arch_add_171_carry_24_, fu_ALU_fu_arch_add_171_carry_25_,
         fu_ALU_fu_arch_add_171_carry_26_, fu_ALU_fu_arch_add_171_carry_27_,
         fu_ALU_fu_arch_add_171_carry_28_, fu_ALU_fu_arch_add_171_carry_29_,
         fu_ALU_fu_arch_add_171_carry_30_, fu_ALU_fu_arch_add_171_carry_31_,
         n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1734, n1735,
         n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1757,
         n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
         n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
         n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
         n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
         n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
         n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
         n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
         n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
         n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
         n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
         n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
         n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
         n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
         n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
         n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
         n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
         n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, fu_LIFTING_n500, fu_LIFTING_n499, fu_LIFTING_n498,
         fu_LIFTING_n497, fu_LIFTING_n496, fu_LIFTING_n495, fu_LIFTING_n494,
         fu_LIFTING_n493, fu_LIFTING_n492, fu_LIFTING_n491, fu_LIFTING_n490,
         fu_LIFTING_n489, fu_LIFTING_n488, fu_LIFTING_n487, fu_LIFTING_n486,
         fu_LIFTING_n485, fu_LIFTING_n484, fu_LIFTING_n483, fu_LIFTING_n482,
         fu_LIFTING_n481, fu_LIFTING_n480, fu_LIFTING_n479, fu_LIFTING_n478,
         fu_LIFTING_n477, fu_LIFTING_n476, fu_LIFTING_n475, fu_LIFTING_n474,
         fu_LIFTING_n473, fu_LIFTING_n472, fu_LIFTING_n471, fu_LIFTING_n470,
         fu_LIFTING_n469, fu_LIFTING_n468, fu_LIFTING_n467, fu_LIFTING_n466,
         fu_LIFTING_n465, fu_LIFTING_n464, fu_LIFTING_n463, fu_LIFTING_n462,
         fu_LIFTING_n461, fu_LIFTING_n460, fu_LIFTING_n459, fu_LIFTING_n458,
         fu_LIFTING_n457, fu_LIFTING_n456, fu_LIFTING_n455, fu_LIFTING_n454,
         fu_LIFTING_n453, fu_LIFTING_n452, fu_LIFTING_n451, fu_LIFTING_n450,
         fu_LIFTING_n449, fu_LIFTING_n448, fu_LIFTING_n447, fu_LIFTING_n446,
         fu_LIFTING_n445, fu_LIFTING_n444, fu_LIFTING_n443, fu_LIFTING_n442,
         fu_LIFTING_n441, fu_LIFTING_n440, fu_LIFTING_n439, fu_LIFTING_n438,
         fu_LIFTING_n437, fu_LIFTING_n436, fu_LIFTING_n435, fu_LIFTING_n434,
         fu_LIFTING_n433, fu_LIFTING_n432, fu_LIFTING_n431, fu_LIFTING_n430,
         fu_LIFTING_n429, fu_LIFTING_n428, fu_LIFTING_n427, fu_LIFTING_n426,
         fu_LIFTING_n425, fu_LIFTING_n424, fu_LIFTING_n423, fu_LIFTING_n422,
         fu_LIFTING_n421, fu_LIFTING_n420, fu_LIFTING_n419, fu_LIFTING_n418,
         fu_LIFTING_n417, fu_LIFTING_n416, fu_LIFTING_n415, fu_LIFTING_n414,
         fu_LIFTING_n413, fu_LIFTING_n412, fu_LIFTING_n411, fu_LIFTING_n410,
         fu_LIFTING_n409, fu_LIFTING_n408, fu_LIFTING_n407, fu_LIFTING_n406,
         fu_LIFTING_n405, fu_LIFTING_n404, fu_LIFTING_n403, fu_LIFTING_n402,
         fu_LIFTING_n401, fu_LIFTING_n400, fu_LIFTING_n399, fu_LIFTING_n398,
         fu_LIFTING_n397, fu_LIFTING_n396, fu_LIFTING_n395, fu_LIFTING_n394,
         fu_LIFTING_n393, fu_LIFTING_n392, fu_LIFTING_n391, fu_LIFTING_n390,
         fu_LIFTING_n389, fu_LIFTING_n388, fu_LIFTING_n387, fu_LIFTING_n386,
         fu_LIFTING_n385, fu_LIFTING_n384, fu_LIFTING_n383, fu_LIFTING_n382,
         fu_LIFTING_n381, fu_LIFTING_n380, fu_LIFTING_n379, fu_LIFTING_n378,
         fu_LIFTING_n377, fu_LIFTING_n376, fu_LIFTING_n375, fu_LIFTING_n374,
         fu_LIFTING_n373, fu_LIFTING_n372, fu_LIFTING_n371, fu_LIFTING_n370,
         fu_LIFTING_n369, fu_LIFTING_n368, fu_LIFTING_n367, fu_LIFTING_n366,
         fu_LIFTING_n365, fu_LIFTING_n364, fu_LIFTING_n363, fu_LIFTING_n362,
         fu_LIFTING_n361, fu_LIFTING_n360, fu_LIFTING_n359, fu_LIFTING_n358,
         fu_LIFTING_n357, fu_LIFTING_n356, fu_LIFTING_n355, fu_LIFTING_n354,
         fu_LIFTING_n353, fu_LIFTING_n352, fu_LIFTING_n351, fu_LIFTING_n350,
         fu_LIFTING_n349, fu_LIFTING_n348, fu_LIFTING_n347, fu_LIFTING_n346,
         fu_LIFTING_n345, fu_LIFTING_n344, fu_LIFTING_n343, fu_LIFTING_n342,
         fu_LIFTING_n341, fu_LIFTING_n340, fu_LIFTING_n339, fu_LIFTING_n338,
         fu_LIFTING_n337, fu_LIFTING_n336, fu_LIFTING_n335, fu_LIFTING_n334,
         fu_LIFTING_n333, fu_LIFTING_n332, fu_LIFTING_n331, fu_LIFTING_n330,
         fu_LIFTING_n329, fu_LIFTING_n328, fu_LIFTING_n327, fu_LIFTING_n326,
         fu_LIFTING_n325, fu_LIFTING_n324, fu_LIFTING_n323, fu_LIFTING_n322,
         fu_LIFTING_n321, fu_LIFTING_n320, fu_LIFTING_n319, fu_LIFTING_n318,
         fu_LIFTING_n317, fu_LIFTING_n316, fu_LIFTING_n315, fu_LIFTING_n314,
         fu_LIFTING_n313, fu_LIFTING_n312, fu_LIFTING_n311, fu_LIFTING_n310,
         fu_LIFTING_n309, fu_LIFTING_n308, fu_LIFTING_n307, fu_LIFTING_n306,
         fu_LIFTING_n305, fu_LIFTING_n304, fu_LIFTING_n303, fu_LIFTING_n302,
         fu_LIFTING_n301, fu_LIFTING_n300, fu_LIFTING_n299, fu_LIFTING_n298,
         fu_LIFTING_n297, fu_LIFTING_n296, fu_LIFTING_n295, fu_LIFTING_n294,
         fu_LIFTING_n293, fu_LIFTING_n292, fu_LIFTING_n291, fu_LIFTING_n290,
         fu_LIFTING_n289, fu_LIFTING_n288, fu_LIFTING_n287, fu_LIFTING_n286,
         fu_LIFTING_n285, fu_LIFTING_n284, fu_LIFTING_n283, fu_LIFTING_n282,
         fu_LIFTING_n281, fu_LIFTING_n280, fu_LIFTING_n279, fu_LIFTING_n278,
         fu_LIFTING_n277, fu_LIFTING_n276, fu_LIFTING_n275, fu_LIFTING_n274,
         fu_LIFTING_n273, fu_LIFTING_n272, fu_LIFTING_n271, fu_LIFTING_n270,
         fu_LIFTING_n269, fu_LIFTING_n268, fu_LIFTING_n267, fu_LIFTING_n266,
         fu_LIFTING_n265, fu_LIFTING_n264, fu_LIFTING_n263, fu_LIFTING_n262,
         fu_LIFTING_n261, fu_LIFTING_n260, fu_LIFTING_n259, fu_LIFTING_n258,
         fu_LIFTING_n257, fu_LIFTING_n256, fu_LIFTING_n255, fu_LIFTING_n254,
         fu_LIFTING_n253, fu_LIFTING_n252, fu_LIFTING_n251, fu_LIFTING_n250,
         fu_LIFTING_n249, fu_LIFTING_n248, fu_LIFTING_n247, fu_LIFTING_n246,
         fu_LIFTING_n245, fu_LIFTING_n244, fu_LIFTING_n243, fu_LIFTING_n242,
         fu_LIFTING_n241, fu_LIFTING_n240, fu_LIFTING_n239, fu_LIFTING_n238,
         fu_LIFTING_n237, fu_LIFTING_n236, fu_LIFTING_n235, fu_LIFTING_n234,
         fu_LIFTING_n233, fu_LIFTING_n231, fu_LIFTING_n135, fu_LIFTING_n134,
         fu_LIFTING_n133, fu_LIFTING_n132, fu_LIFTING_n131, fu_LIFTING_n130,
         fu_LIFTING_n129, fu_LIFTING_n128, fu_LIFTING_n127, fu_LIFTING_n126,
         fu_LIFTING_n125, fu_LIFTING_n124, fu_LIFTING_n123, fu_LIFTING_n122,
         fu_LIFTING_n121, fu_LIFTING_n120, fu_LIFTING_n119, fu_LIFTING_n118,
         fu_LIFTING_n117, fu_LIFTING_n116, fu_LIFTING_n115, fu_LIFTING_n114,
         fu_LIFTING_n113, fu_LIFTING_n112, fu_LIFTING_n111, fu_LIFTING_n110,
         fu_LIFTING_n109, fu_LIFTING_n108, fu_LIFTING_n106, fu_LIFTING_n105,
         fu_LIFTING_n104, fu_LIFTING_n103, fu_LIFTING_n102, fu_LIFTING_n101,
         fu_LIFTING_n100, fu_LIFTING_n99, fu_LIFTING_n98, fu_LIFTING_n97,
         fu_LIFTING_n96, fu_LIFTING_n95, fu_LIFTING_n94, fu_LIFTING_n93,
         fu_LIFTING_n92, fu_LIFTING_n91, fu_LIFTING_n90, fu_LIFTING_n89,
         fu_LIFTING_n88, fu_LIFTING_n87, fu_LIFTING_n85, fu_LIFTING_n84,
         fu_LIFTING_n83, fu_LIFTING_n82, fu_LIFTING_n81, fu_LIFTING_n80,
         fu_LIFTING_n79, fu_LIFTING_n78, fu_LIFTING_n77, fu_LIFTING_n76,
         fu_LIFTING_n73, fu_LIFTING_n71, fu_LIFTING_n70, fu_LIFTING_n69,
         fu_LIFTING_n68, fu_LIFTING_n67, fu_LIFTING_n66, fu_LIFTING_n65,
         fu_LIFTING_n64, fu_LIFTING_n63, fu_LIFTING_n62, fu_LIFTING_n61,
         fu_LIFTING_n60, fu_LIFTING_n59, fu_LIFTING_n58, fu_LIFTING_n57,
         fu_LIFTING_n56, fu_LIFTING_n55, fu_LIFTING_n54, fu_LIFTING_n53,
         fu_LIFTING_n52, fu_LIFTING_n51, fu_LIFTING_n50, fu_LIFTING_n49,
         fu_LIFTING_n48, fu_LIFTING_n47, fu_LIFTING_n46, fu_LIFTING_n45,
         fu_LIFTING_n44, fu_LIFTING_n43, fu_LIFTING_n42, fu_LIFTING_n41,
         fu_LIFTING_n40, fu_LIFTING_n39, fu_LIFTING_n37, fu_LIFTING_n36,
         fu_LIFTING_n3, fu_LIFTING_n2, fu_LIFTING_n1,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n1,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n2,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n3,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n4,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n5,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n6,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n7,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n8,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n9,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n10,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n11,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n12,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n13,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n14,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n15,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n16,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n17,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n18,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n19,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n20,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n21,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n22,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n23,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n24,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n25,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n26,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n27,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n28,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n29,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n30,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n31,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n32,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n39,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n40,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n41,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n42,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n43,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n44,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n45,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n46,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n47,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n48,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n49,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n50,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n51,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n52,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n53,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n54,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n55,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n56,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n57,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n58,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n59,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n60,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n61,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n62,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n63,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n64,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n65,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n66,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n67,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n68,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n69,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n70,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n71,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_n72,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_0_,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_1_,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_2_,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_3_,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_4_,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_5_,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_6_,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_7_,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_8_,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_9_,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_10_,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_11_,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_12_,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_13_,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_14_,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_15_,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_16_,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_17_,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_18_,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_19_,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_20_,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_21_,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_22_,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_23_,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_24_,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_25_,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_26_,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_27_,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_28_,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_29_,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_30_,
         fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_31_,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n2,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n3,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n4,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n5,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n6,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n7,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n8,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n9,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n10,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n11,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n12,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n13,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n14,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n15,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n16,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n17,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n18,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n19,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n20,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n21,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n22,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n23,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n24,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n25,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n36,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n37,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n38,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n39,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n40,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n41,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n42,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n43,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n44,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n45,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n46,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n47,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n48,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n49,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n50,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n51,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n52,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n53,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n54,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n55,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n56,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n57,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n58,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n59,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n60,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n61,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n62,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n63,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n64,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n65,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n66,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n67,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n68,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n69,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n70,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n71,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n72,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n73,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n74,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n75,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n76,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n77,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n78,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n79,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n80,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n81,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n82,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n83,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n84,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n85,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n86,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n87,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n88,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n89,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n90,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n91,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n92,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n93,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n94,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n95,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n96,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n97,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n98,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n99,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n100,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n101,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n102,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n103,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n104,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n105,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n106,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n107,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n108,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n109,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n110,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n111,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n112,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n113,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n114,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n115,
         fu_LIFTING_mult_75_DP_OP_278_6650_1_n116,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n2,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n3,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n4,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n5,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n6,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n7,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n8,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n9,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n10,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n11,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n12,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n13,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n14,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n15,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n16,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n17,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n18,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n19,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n20,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n21,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n22,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n23,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n24,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n25,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n29,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n30,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n31,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n32,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n33,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n34,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n35,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n36,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n37,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n38,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n39,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n40,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n41,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n42,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n43,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n44,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n45,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n46,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n47,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n48,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n49,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n50,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n51,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n52,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n53,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n54,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n55,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n56,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n57,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n58,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n59,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n60,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n61,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n62,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n63,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n64,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n65,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n66,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n67,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n68,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n69,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n70,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n71,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n72,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n73,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n74,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n75,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n76,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n77,
         fu_LIFTING_mult_79_DP_OP_279_6650_2_n78,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n2,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n3,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n4,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n5,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n6,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n7,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n8,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n9,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n10,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n11,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n12,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n13,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n14,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n15,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n16,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n17,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n18,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n19,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n20,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n21,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n22,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n23,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n24,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n25,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n31,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n32,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n33,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n34,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n35,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n36,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n37,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n38,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n39,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n40,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n41,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n42,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n43,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n44,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n45,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n46,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n47,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n48,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n49,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n50,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n51,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n52,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n53,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n54,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n55,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n56,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n57,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n58,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n59,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n60,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n61,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n62,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n63,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n64,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n65,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n66,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n67,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n68,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n69,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n70,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n71,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n72,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n73,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n74,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n75,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n76,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n77,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n78,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n79,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n80,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n81,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n82,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n83,
         fu_LIFTING_mult_84_DP_OP_276_6650_3_n84,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n2,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n3,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n4,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n5,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n6,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n7,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n8,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n9,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n10,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n11,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n12,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n13,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n14,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n15,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n16,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n17,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n18,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n19,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n20,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n21,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n22,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n23,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n24,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n25,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n30,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n31,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n32,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n33,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n34,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n35,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n36,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n37,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n38,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n39,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n40,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n41,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n42,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n43,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n44,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n45,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n46,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n47,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n48,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n49,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n50,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n51,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n52,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n53,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n54,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n55,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n56,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n57,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n58,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n59,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n60,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n61,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n62,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n63,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n64,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n65,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n66,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n67,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n68,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n69,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n70,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n71,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n72,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n73,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n74,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n75,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n76,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n77,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n78,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n79,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n80,
         fu_LIFTING_mult_88_DP_OP_277_6650_4_n81,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n2,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n3,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n4,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n5,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n6,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n7,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n8,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n9,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n10,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n11,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n12,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n13,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n14,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n15,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n16,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n17,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n18,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n19,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n20,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n21,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n22,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n23,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n24,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n25,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n33,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n34,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n35,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n36,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n37,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n38,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n39,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n40,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n41,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n42,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n43,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n44,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n45,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n46,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n47,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n48,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n49,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n50,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n51,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n52,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n53,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n54,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n55,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n56,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n57,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n58,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n59,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n60,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n61,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n62,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n63,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n64,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n65,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n66,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n67,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n68,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n69,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n70,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n71,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n72,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n73,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n74,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n75,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n76,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n77,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n78,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n79,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n80,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n81,
         fu_LIFTING_mult_92_DP_OP_280_6650_5_n82,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n2,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n3,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n4,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n5,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n6,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n7,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n8,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n9,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n10,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n11,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n12,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n13,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n14,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n15,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n16,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n17,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n18,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n19,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n20,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n21,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n22,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n23,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n24,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n25,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n33,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n34,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n35,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n36,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n37,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n38,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n39,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n40,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n41,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n42,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n43,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n44,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n45,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n46,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n47,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n48,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n49,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n50,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n51,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n52,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n53,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n54,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n55,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n56,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n57,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n58,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n59,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n60,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n61,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n62,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n63,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n64,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n65,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n66,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n67,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n68,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n69,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n70,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n71,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n72,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n73,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n74,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n75,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n76,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n77,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n78,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n79,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n80,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n82,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n83,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n86,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n88,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n89,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n90,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n91,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n92,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n94,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n95,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n97,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n99,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n100,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n102,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n103,
         fu_LIFTING_mult_96_DP_OP_281_6650_6_n104, fu_LIFTING_n107,
         fu_LIFTING_n75, fu_LIFTING_n74, fu_LIFTING_n72, fu_LIFTING_N993,
         fu_LIFTING_N961, fu_LIFTING_N929, fu_LIFTING_N703, fu_LIFTING_N702,
         fu_LIFTING_N701, fu_LIFTING_N700, fu_LIFTING_N699, fu_LIFTING_N698,
         fu_LIFTING_N697, fu_LIFTING_N696, fu_LIFTING_N695, fu_LIFTING_N694,
         fu_LIFTING_N693, fu_LIFTING_N692, fu_LIFTING_N691, fu_LIFTING_N690,
         fu_LIFTING_N689, fu_LIFTING_N688, fu_LIFTING_N687, fu_LIFTING_N686,
         fu_LIFTING_N685, fu_LIFTING_N684, fu_LIFTING_N683, fu_LIFTING_N682,
         fu_LIFTING_N681, fu_LIFTING_N680, fu_LIFTING_N679, fu_LIFTING_N678,
         fu_LIFTING_N677, fu_LIFTING_N676, fu_LIFTING_N675, fu_LIFTING_N674,
         fu_LIFTING_N673, fu_LIFTING_N672, fu_LIFTING_N671, fu_LIFTING_N670,
         fu_LIFTING_N669, fu_LIFTING_N668, fu_LIFTING_N667, fu_LIFTING_N666,
         fu_LIFTING_N665, fu_LIFTING_N664, fu_LIFTING_N663, fu_LIFTING_N662,
         fu_LIFTING_N661, fu_LIFTING_N660, fu_LIFTING_N659, fu_LIFTING_N658,
         fu_LIFTING_N657, fu_LIFTING_N656, fu_LIFTING_N655, fu_LIFTING_N654,
         fu_LIFTING_N653, fu_LIFTING_N652, fu_LIFTING_N651, fu_LIFTING_N650,
         fu_LIFTING_N649, fu_LIFTING_N648, fu_LIFTING_N647, fu_LIFTING_N646,
         fu_LIFTING_N645, fu_LIFTING_N644, fu_LIFTING_N551, fu_LIFTING_N550,
         fu_LIFTING_N549, fu_LIFTING_N548, fu_LIFTING_N547, fu_LIFTING_N546,
         fu_LIFTING_N545, fu_LIFTING_N544, fu_LIFTING_N543, fu_LIFTING_N542,
         fu_LIFTING_N541, fu_LIFTING_N540, fu_LIFTING_N539, fu_LIFTING_N538,
         fu_LIFTING_N537, fu_LIFTING_N536, fu_LIFTING_N535, fu_LIFTING_N534,
         fu_LIFTING_N533, fu_LIFTING_N532, fu_LIFTING_N531, fu_LIFTING_N530,
         fu_LIFTING_N529, fu_LIFTING_N528, fu_LIFTING_N431, fu_LIFTING_N430,
         fu_LIFTING_N429, fu_LIFTING_N428, fu_LIFTING_N427, fu_LIFTING_N426,
         fu_LIFTING_N425, fu_LIFTING_N424, fu_LIFTING_N423, fu_LIFTING_N422,
         fu_LIFTING_N421, fu_LIFTING_N420, fu_LIFTING_N419, fu_LIFTING_N418,
         fu_LIFTING_N417, fu_LIFTING_N416, fu_LIFTING_N415, fu_LIFTING_N414,
         fu_LIFTING_N413, fu_LIFTING_N412, fu_LIFTING_N411, fu_LIFTING_N410,
         fu_LIFTING_N409, fu_LIFTING_N408, fu_LIFTING_N311, fu_LIFTING_N310,
         fu_LIFTING_N309, fu_LIFTING_N308, fu_LIFTING_N307, fu_LIFTING_N306,
         fu_LIFTING_N305, fu_LIFTING_N304, fu_LIFTING_N303, fu_LIFTING_N302,
         fu_LIFTING_N301, fu_LIFTING_N300, fu_LIFTING_N299, fu_LIFTING_N298,
         fu_LIFTING_N297, fu_LIFTING_N296, fu_LIFTING_N295, fu_LIFTING_N294,
         fu_LIFTING_N293, fu_LIFTING_N292, fu_LIFTING_N291, fu_LIFTING_N290,
         fu_LIFTING_N289, fu_LIFTING_N288, fu_LIFTING_N191, fu_LIFTING_N190,
         fu_LIFTING_N189, fu_LIFTING_N188, fu_LIFTING_N187, fu_LIFTING_N186,
         fu_LIFTING_N185, fu_LIFTING_N184, fu_LIFTING_N183, fu_LIFTING_N182,
         fu_LIFTING_N181, fu_LIFTING_N180, fu_LIFTING_N179, fu_LIFTING_N178,
         fu_LIFTING_N177, fu_LIFTING_N176, fu_LIFTING_N175, fu_LIFTING_N174,
         fu_LIFTING_N173, fu_LIFTING_N172, fu_LIFTING_N171, fu_LIFTING_N170,
         fu_LIFTING_N169, fu_LIFTING_N168, fu_LIFTING_reg_out_tmp_0_,
         fu_LIFTING_reg_out_tmp_1_, fu_LIFTING_reg_out_tmp_2_,
         fu_LIFTING_reg_out_tmp_3_, fu_LIFTING_reg_out_tmp_4_,
         fu_LIFTING_reg_out_tmp_5_, fu_LIFTING_reg_out_tmp_6_,
         fu_LIFTING_reg_out_tmp_7_, fu_LIFTING_reg_out_tmp_8_,
         fu_LIFTING_reg_out_tmp_9_, fu_LIFTING_reg_out_tmp_10_,
         fu_LIFTING_reg_out_tmp_11_, fu_LIFTING_reg_out_tmp_12_,
         fu_LIFTING_reg_out_tmp_13_, fu_LIFTING_reg_out_tmp_14_,
         fu_LIFTING_reg_out_tmp_15_, fu_LIFTING_reg_out_tmp_16_,
         fu_LIFTING_reg_out_tmp_17_, fu_LIFTING_reg_out_tmp_18_,
         fu_LIFTING_reg_out_tmp_19_, fu_LIFTING_reg_out_tmp_20_,
         fu_LIFTING_reg_out_tmp_21_, fu_LIFTING_reg_out_tmp_22_,
         fu_LIFTING_reg_out_tmp_23_, fu_LIFTING_reg_out_tmp_24_,
         fu_LIFTING_reg_out_tmp_25_, fu_LIFTING_reg_out_tmp_26_,
         fu_LIFTING_reg_out_tmp_27_, fu_LIFTING_reg_out_tmp_28_,
         fu_LIFTING_reg_out_tmp_29_, fu_LIFTING_reg_out_tmp_30_,
         fu_LIFTING_reg_out_tmp_31_, fu_LIFTING_N99, fu_LIFTING_N98,
         fu_LIFTING_N97, fu_LIFTING_N96, fu_LIFTING_N95, fu_LIFTING_N94,
         fu_LIFTING_N93, fu_LIFTING_N92, fu_LIFTING_N91, fu_LIFTING_N90,
         fu_LIFTING_N89, fu_LIFTING_N88, fu_LIFTING_N87, fu_LIFTING_N86,
         fu_LIFTING_N85, fu_LIFTING_N84, fu_LIFTING_N83, fu_LIFTING_N82,
         fu_LIFTING_N81, fu_LIFTING_N80, fu_LIFTING_N79, fu_LIFTING_N78,
         fu_LIFTING_N77, fu_LIFTING_N76, fu_LIFTING_N75, fu_LIFTING_N74,
         fu_LIFTING_N73, fu_LIFTING_N72, fu_LIFTING_N71, fu_LIFTING_N70,
         fu_LIFTING_N69, fu_LIFTING_N68, fu_LIFTING_N67, fu_LIFTING_N66,
         fu_LIFTING_N65, fu_LIFTING_N64, fu_LIFTING_N63, fu_LIFTING_N62,
         fu_LIFTING_N61, fu_LIFTING_N60, fu_LIFTING_N59, fu_LIFTING_N58,
         fu_LIFTING_N57, fu_LIFTING_N56, fu_LIFTING_N55, fu_LIFTING_N54,
         fu_LIFTING_N53, fu_LIFTING_N52, fu_LIFTING_N51, fu_LIFTING_N50,
         fu_LIFTING_N49, fu_LIFTING_N48, fu_LIFTING_reg_x1_0_,
         fu_LIFTING_reg_x1_1_, fu_LIFTING_reg_x1_2_, fu_LIFTING_reg_x1_3_,
         fu_LIFTING_reg_x1_4_, fu_LIFTING_reg_x1_5_, fu_LIFTING_reg_x1_6_,
         fu_LIFTING_reg_x1_7_, fu_LIFTING_reg_x1_8_, fu_LIFTING_reg_x1_9_,
         fu_LIFTING_reg_x1_10_, fu_LIFTING_reg_x1_11_, fu_LIFTING_reg_x1_12_,
         fu_LIFTING_reg_x1_13_, fu_LIFTING_reg_x1_14_, fu_LIFTING_reg_x1_15_,
         fu_LIFTING_reg_x1_16_, fu_LIFTING_reg_x1_17_, fu_LIFTING_reg_x1_18_,
         fu_LIFTING_reg_x1_19_, fu_LIFTING_reg_x1_20_, fu_LIFTING_reg_x1_21_,
         fu_LIFTING_reg_x1_22_, fu_LIFTING_reg_x1_23_, fu_LIFTING_reg_x1_24_,
         fu_LIFTING_reg_x1_25_, fu_LIFTING_reg_x1_26_, fu_LIFTING_reg_x1_27_,
         fu_LIFTING_reg_x1_28_, fu_LIFTING_reg_x1_29_, fu_LIFTING_reg_x1_30_,
         fu_LIFTING_reg_x1_31_, fu_LIFTING_reg_x2_0_, fu_LIFTING_reg_x2_1_,
         fu_LIFTING_reg_x2_2_, fu_LIFTING_reg_x2_3_, fu_LIFTING_reg_x2_4_,
         fu_LIFTING_reg_x2_5_, fu_LIFTING_reg_x2_6_, fu_LIFTING_reg_x2_7_,
         fu_LIFTING_reg_x2_8_, fu_LIFTING_reg_x2_9_, fu_LIFTING_reg_x2_10_,
         fu_LIFTING_reg_x2_11_, fu_LIFTING_reg_x2_12_, fu_LIFTING_reg_x2_13_,
         fu_LIFTING_reg_x2_14_, fu_LIFTING_reg_x2_15_, fu_LIFTING_reg_x2_16_,
         fu_LIFTING_reg_x2_17_, fu_LIFTING_reg_x2_18_, fu_LIFTING_reg_x2_19_,
         fu_LIFTING_reg_x2_20_, fu_LIFTING_reg_x2_21_, fu_LIFTING_reg_x2_22_,
         fu_LIFTING_reg_x2_23_, fu_LIFTING_reg_x2_24_, fu_LIFTING_reg_x2_25_,
         fu_LIFTING_reg_x2_26_, fu_LIFTING_reg_x2_27_, fu_LIFTING_reg_x2_28_,
         fu_LIFTING_reg_x2_29_, fu_LIFTING_reg_x2_30_, fu_LIFTING_reg_x2_31_;
  wire   [14:0] ic_socket_gcu_o1_data0_wire;
  wire   [41:0] inst_decoder_instructionword_wire;
  wire   [31:0] ic_simm_B1_wire;
  wire   [2:0] fu_LSU_t1opcode_wire;
  wire   [3:0] fu_ALU_t1opcode_wire;
  wire   [2:0] fu_LIFTING_t1opcode_wire;
  wire   [2:0] rf_RF_t1opcode_wire;
  wire   [2:0] rf_RF_r1opcode_wire;
  wire   [31:0] ic_socket_lsu_o1_data0_wire;
  wire   [31:0] ic_socket_ALU_o1_data0_wire;
  wire   [31:0] ic_socket_LIFTING_o1_data0_wire;
  wire   [31:0] rf_RF_t1data_wire;
  wire   [0:31] fu_ALU_o1reg;
  wire   [0:3] fu_ALU_opc1reg;
  wire   [2:31] fu_ALU_t1reg;
  assign imem_en_x = 1'b0;

  OAI211X4 U1133 ( .A0(inst_decoder_instructionword_wire[40]), .A1(n593), .B0(
        n2210), .C0(n594), .Y(n571) );
  DFFRQX4 fu_ALU_o1reg_reg_11_ ( .D(n843), .CK(clk), .RN(rstx), .Q(
        fu_ALU_o1reg[11]) );
  OAI22X1 fu_ALU_fu_arch_U500 ( .A0(n2093), .A1(n1738), .B0(n1776), .B1(n1773), 
        .Y(fu_ALU_fu_arch_n691) );
  OAI21X1 fu_ALU_fu_arch_U235 ( .A0(n2139), .A1(n2195), .B0(
        fu_ALU_fu_arch_n475), .Y(fu_ALU_fu_arch_n473) );
  AOI221X2 fu_ALU_fu_arch_U150 ( .A0(n2188), .A1(n2128), .B0(
        fu_ALU_fu_arch_n175), .B1(n1765), .C0(n2190), .Y(fu_ALU_fu_arch_n356)
         );
  AOI31X1 fu_ALU_fu_arch_U143 ( .A0(fu_ALU_fu_arch_n348), .A1(
        fu_ALU_fu_arch_n349), .A2(fu_ALU_fu_arch_n350), .B0(
        fu_ALU_fu_arch_n308), .Y(fu_ALU_fu_arch_n341) );
  AOI221X2 fu_ALU_fu_arch_U163 ( .A0(n2188), .A1(n2130), .B0(
        fu_ALU_fu_arch_n175), .B1(n1747), .C0(n2190), .Y(fu_ALU_fu_arch_n376)
         );
  OAI21X1 fu_ALU_fu_arch_U287 ( .A0(n2145), .A1(n2195), .B0(
        fu_ALU_fu_arch_n529), .Y(fu_ALU_fu_arch_n528) );
  AOI221X2 fu_ALU_fu_arch_U401 ( .A0(n1762), .A1(n1767), .B0(n2188), .B1(n2154), .C0(n2190), .Y(fu_ALU_fu_arch_n629) );
  AOI31X1 fu_ALU_fu_arch_U422 ( .A0(n2179), .A1(n2155), .A2(
        fu_ALU_fu_arch_n175), .B0(fu_ALU_fu_arch_n128), .Y(fu_ALU_fu_arch_n650) );
  AOI31X1 fu_ALU_fu_arch_U438 ( .A0(n2156), .A1(fu_ALU_fu_arch_n621), .A2(
        n1762), .B0(fu_ALU_fu_arch_n128), .Y(fu_ALU_fu_arch_n663) );
  OAI22X1 fu_ALU_fu_arch_U488 ( .A0(fu_ALU_fu_arch_n372), .A1(
        fu_ALU_fu_arch_n212), .B0(fu_ALU_fu_arch_n155), .B1(
        fu_ALU_fu_arch_n138), .Y(fu_ALU_fu_arch_n678) );
  AOI31X1 fu_ALU_fu_arch_U505 ( .A0(n2160), .A1(n2159), .A2(n1762), .B0(
        fu_ALU_fu_arch_n128), .Y(fu_ALU_fu_arch_n698) );
  AOI31X1 fu_ALU_fu_arch_U550 ( .A0(n2162), .A1(n1772), .A2(
        fu_ALU_fu_arch_n175), .B0(fu_ALU_fu_arch_n128), .Y(fu_ALU_fu_arch_n721) );
  AOI31X1 fu_ALU_fu_arch_U16 ( .A0(n1762), .A1(n2163), .A2(n1778), .B0(
        fu_ALU_fu_arch_n128), .Y(fu_ALU_fu_arch_n127) );
  AOI221X2 fu_ALU_fu_arch_U14 ( .A0(n2188), .A1(n2163), .B0(n1762), .B1(n1745), 
        .C0(n2190), .Y(fu_ALU_fu_arch_n119) );
  OAI22X1 fu_ALU_fu_arch_U40 ( .A0(fu_ALU_fu_arch_n154), .A1(
        fu_ALU_fu_arch_n132), .B0(fu_ALU_fu_arch_n155), .B1(
        fu_ALU_fu_arch_n134), .Y(fu_ALU_fu_arch_n144) );
  AOI31X1 fu_ALU_fu_arch_U35 ( .A0(n1762), .A1(n2165), .A2(n2164), .B0(
        fu_ALU_fu_arch_n128), .Y(fu_ALU_fu_arch_n152) );
  AOI221X2 fu_ALU_fu_arch_U33 ( .A0(n2188), .A1(n2165), .B0(n1762), .B1(n1742), 
        .C0(n2190), .Y(fu_ALU_fu_arch_n148) );
  AOI221X2 fu_ALU_fu_arch_U47 ( .A0(n1762), .A1(n1766), .B0(n2188), .B1(n2167), 
        .C0(n2190), .Y(fu_ALU_fu_arch_n172) );
  AOI221X2 fu_ALU_fu_arch_U55 ( .A0(n1762), .A1(n1741), .B0(n2099), .B1(n2169), 
        .C0(n2190), .Y(fu_ALU_fu_arch_n186) );
  AOI221X2 fu_ALU_fu_arch_U66 ( .A0(n2188), .A1(fu_ALU_t1reg[5]), .B0(n1762), 
        .B1(n2039), .C0(n2190), .Y(fu_ALU_fu_arch_n205) );
  OAI22X1 fu_ALU_fu_arch_U65 ( .A0(fu_ALU_fu_arch_n204), .A1(
        fu_ALU_fu_arch_n108), .B0(fu_ALU_fu_arch_n205), .B1(n1754), .Y(
        fu_ALU_fu_arch_n203) );
  AOI221X2 fu_ALU_fu_arch_U76 ( .A0(fu_ALU_fu_arch_n175), .A1(
        fu_ALU_fu_arch_n220), .B0(n2188), .B1(n2172), .C0(n2190), .Y(
        fu_ALU_fu_arch_n221) );
  AOI221X2 fu_ALU_fu_arch_U85 ( .A0(n1762), .A1(n1768), .B0(n2188), .B1(n2174), 
        .C0(n2190), .Y(fu_ALU_fu_arch_n236) );
  AOI221X2 fu_ALU_fu_arch_U136 ( .A0(n1762), .A1(fu_ALU_fu_arch_n335), .B0(
        n2099), .B1(n2176), .C0(n2190), .Y(fu_ALU_fu_arch_n331) );
  OAI22X1 fu_ALU_fu_arch_U130 ( .A0(n2107), .A1(n1754), .B0(n1776), .B1(n1773), 
        .Y(fu_ALU_fu_arch_n322) );
  OAI22X1 fu_ALU_fu_arch_U129 ( .A0(n1769), .A1(n2171), .B0(n2199), .B1(n2175), 
        .Y(fu_ALU_fu_arch_n323) );
  OAI21X1 fu_ALU_fu_arch_U128 ( .A0(fu_ALU_fu_arch_n322), .A1(
        fu_ALU_fu_arch_n323), .B0(fu_ALU_fu_arch_n249), .Y(fu_ALU_fu_arch_n320) );
  AOI221X2 fu_ALU_fu_arch_U313 ( .A0(n2099), .A1(fu_ALU_fu_arch_sub_200_A_1_), 
        .B0(fu_ALU_fu_arch_n175), .B1(n1770), .C0(n2190), .Y(
        fu_ALU_fu_arch_n556) );
  NOR2X8 fu_ALU_fu_arch_U706 ( .A(fu_ALU_fu_arch_n746), .B(fu_ALU_fu_arch_n761), .Y(fu_ALU_fu_arch_n274) );
  AOI211X4 fu_ALU_fu_arch_U663 ( .A0(n2136), .A1(n2198), .B0(
        fu_ALU_fu_arch_n310), .C0(fu_ALU_fu_arch_n764), .Y(fu_ALU_fu_arch_n535) );
  AOI21X1 fu_ALU_fu_arch_U218 ( .A0(n2188), .A1(n2137), .B0(n2190), .Y(
        fu_ALU_fu_arch_n452) );
  OAI21X1 fu_ALU_fu_arch_U217 ( .A0(n2137), .A1(n2196), .B0(
        fu_ALU_fu_arch_n452), .Y(fu_ALU_fu_arch_n450) );
  OR3X2 fu_ALU_fu_arch_U610 ( .A(fu_ALU_fu_arch_n744), .B(fu_ALU_fu_arch_n745), 
        .C(fu_ALU_opc1reg[0]), .Y(fu_ALU_fu_arch_n631) );
  OAI211X4 fu_ALU_fu_arch_U530 ( .A0(n1764), .A1(n2199), .B0(
        fu_ALU_fu_arch_n707), .C0(fu_ALU_fu_arch_n708), .Y(fu_ALU_fu_arch_n481) );
  AOI22X1 fu_ALU_fu_arch_U173 ( .A0(n2201), .A1(fu_ALU_o1reg[25]), .B0(n2200), 
        .B1(n2132), .Y(fu_ALU_fu_arch_n392) );
  AOI22X1 fu_ALU_fu_arch_U186 ( .A0(n2201), .A1(fu_ALU_o1reg[24]), .B0(n2200), 
        .B1(fu_ALU_o1reg[25]), .Y(fu_ALU_fu_arch_n411) );
  NOR2X1 fu_ALU_fu_arch_U122 ( .A(n2199), .B(n2125), .Y(fu_ALU_fu_arch_n311)
         );
  AOI221X2 U177 ( .A0(ic_simm_B1_wire[23]), .A1(ic_simm_cntrl_B1_wire_0_), 
        .B0(n2219), .B1(rf_RF_reg_0__23_), .C0(n148), .Y(n146) );
  OAI211X4 fu_ALU_fu_arch_U542 ( .A0(n1763), .A1(n2093), .B0(
        fu_ALU_fu_arch_n713), .C0(fu_ALU_fu_arch_n714), .Y(fu_ALU_fu_arch_n482) );
  AOI21X1 fu_ALU_fu_arch_U236 ( .A0(n2188), .A1(n2139), .B0(n2190), .Y(
        fu_ALU_fu_arch_n475) );
  OAI21X6 fu_ALU_fu_arch_U473 ( .A0(n1770), .A1(n1774), .B0(
        fu_ALU_fu_arch_n675), .Y(fu_ALU_fu_arch_n438) );
  OAI21X1 fu_ALU_fu_arch_U441 ( .A0(n1798), .A1(fu_ALU_fu_arch_n544), .B0(
        fu_ALU_fu_arch_n665), .Y(fu_ALU_fu_arch_n664) );
  AOI221X2 U65 ( .A0(ic_simm_B1_wire[28]), .A1(n2258), .B0(n2219), .B1(
        rf_RF_reg_0__28_), .C0(n82), .Y(n80) );
  AOI31X1 fu_ALU_fu_arch_U156 ( .A0(fu_ALU_fu_arch_n369), .A1(
        fu_ALU_fu_arch_n370), .A2(fu_ALU_fu_arch_n371), .B0(
        fu_ALU_fu_arch_n308), .Y(fu_ALU_fu_arch_n362) );
  AND4X4 fu_ALU_fu_arch_U460 ( .A(fu_ALU_fu_arch_n422), .B(fu_ALU_fu_arch_n670), .C(fu_ALU_fu_arch_n393), .D(fu_ALU_fu_arch_n467), .Y(fu_ALU_fu_arch_n135) );
  AOI22X1 U242 ( .A0(n2217), .A1(rf_RF_reg_3__20_), .B0(n2215), .B1(
        rf_RF_reg_1__20_), .Y(n188) );
  AOI221X2 U240 ( .A0(ic_simm_B1_wire[20]), .A1(n2258), .B0(n2219), .B1(
        rf_RF_reg_0__20_), .C0(n185), .Y(n183) );
  AOI21X1 fu_ALU_fu_arch_U288 ( .A0(n2188), .A1(n2145), .B0(n2190), .Y(
        fu_ALU_fu_arch_n529) );
  AOI22X1 fu_ALU_fu_arch_U541 ( .A0(n2198), .A1(fu_ALU_fu_arch_sub_200_B_19_), 
        .B0(n2201), .B1(fu_ALU_o1reg[21]), .Y(fu_ALU_fu_arch_n711) );
  OAI211X4 fu_ALU_fu_arch_U539 ( .A0(n2140), .A1(n2109), .B0(
        fu_ALU_fu_arch_n711), .C0(fu_ALU_fu_arch_n712), .Y(fu_ALU_fu_arch_n167) );
  OR2X4 fu_ALU_fu_arch_U387 ( .A(fu_ALU_fu_arch_n388), .B(n2106), .Y(
        fu_ALU_fu_arch_n563) );
  OAI22X1 fu_ALU_fu_arch_U318 ( .A0(fu_ALU_fu_arch_n234), .A1(
        fu_ALU_fu_arch_n563), .B0(fu_ALU_fu_arch_n564), .B1(n2146), .Y(
        fu_ALU_fu_arch_n562) );
  AOI22X1 U285 ( .A0(n2217), .A1(rf_RF_reg_3__18_), .B0(n2216), .B1(
        rf_RF_reg_1__18_), .Y(n214) );
  OAI22X1 fu_ALU_fu_arch_U338 ( .A0(n1802), .A1(fu_ALU_fu_arch_n563), .B0(
        fu_ALU_fu_arch_n581), .B1(n2148), .Y(fu_ALU_fu_arch_n579) );
  OAI22X1 fu_ALU_fu_arch_U356 ( .A0(n1798), .A1(fu_ALU_fu_arch_n563), .B0(
        n1864), .B1(fu_ALU_fu_arch_n522), .Y(fu_ALU_fu_arch_n596) );
  AOI221X2 U330 ( .A0(ic_simm_B1_wire[16]), .A1(n2258), .B0(n2219), .B1(
        rf_RF_reg_0__16_), .C0(n244), .Y(n242) );
  OAI211X4 fu_ALU_fu_arch_U681 ( .A0(n1776), .A1(fu_ALU_fu_arch_n522), .B0(
        fu_ALU_fu_arch_n766), .C0(fu_ALU_fu_arch_n524), .Y(fu_ALU_fu_arch_n224) );
  AOI22X1 U354 ( .A0(n2217), .A1(rf_RF_reg_3__15_), .B0(n2216), .B1(
        rf_RF_reg_1__15_), .Y(n259) );
  AOI22X1 fu_ALU_fu_arch_U537 ( .A0(n2198), .A1(n2153), .B0(n2202), .B1(
        fu_ALU_fu_arch_sub_200_B_18_), .Y(fu_ALU_fu_arch_n709) );
  NOR2X6 fu_ALU_fu_arch_U483 ( .A(n2106), .B(fu_ALU_fu_arch_n118), .Y(
        fu_ALU_fu_arch_n636) );
  OAI22X1 fu_ALU_fu_arch_U415 ( .A0(fu_ALU_fu_arch_n291), .A1(
        fu_ALU_fu_arch_n212), .B0(fu_ALU_fu_arch_n645), .B1(n2155), .Y(
        fu_ALU_fu_arch_n644) );
  AOI22X1 fu_ALU_fu_arch_U481 ( .A0(n2158), .A1(n2189), .B0(n2196), .B1(n1744), 
        .Y(fu_ALU_fu_arch_n683) );
  OAI21X1 fu_ALU_fu_arch_U480 ( .A0(n2190), .A1(fu_ALU_fu_arch_n683), .B0(
        fu_ALU_o1reg[12]), .Y(fu_ALU_fu_arch_n682) );
  AOI22X1 fu_ALU_fu_arch_U595 ( .A0(n2201), .A1(n2157), .B0(n2200), .B1(
        fu_ALU_fu_arch_sub_200_B_11_), .Y(fu_ALU_fu_arch_n734) );
  NAND2X1 fu_ALU_fu_arch_U305 ( .A(n2197), .B(fu_ALU_fu_arch_sub_200_B_9_), 
        .Y(fu_ALU_fu_arch_n545) );
  OAI22X1 fu_ALU_fu_arch_U20 ( .A0(fu_ALU_fu_arch_n135), .A1(
        fu_ALU_fu_arch_n136), .B0(fu_ALU_fu_arch_n137), .B1(
        fu_ALU_fu_arch_n138), .Y(fu_ALU_fu_arch_n113) );
  OAI22X1 fu_ALU_fu_arch_U13 ( .A0(fu_ALU_fu_arch_n117), .A1(
        fu_ALU_fu_arch_n118), .B0(fu_ALU_fu_arch_n119), .B1(n1778), .Y(
        fu_ALU_fu_arch_n116) );
  OAI22X1 fu_ALU_fu_arch_U41 ( .A0(fu_ALU_fu_arch_n156), .A1(
        fu_ALU_fu_arch_n136), .B0(fu_ALU_fu_arch_n157), .B1(
        fu_ALU_fu_arch_n138), .Y(fu_ALU_fu_arch_n143) );
  OAI22X1 fu_ALU_fu_arch_U32 ( .A0(fu_ALU_fu_arch_n147), .A1(
        fu_ALU_fu_arch_n118), .B0(fu_ALU_fu_arch_n148), .B1(n2164), .Y(
        fu_ALU_fu_arch_n146) );
  NAND4X8 U532 ( .A(n337), .B(n338), .C(n339), .D(n340), .Y(
        rf_RF_t1data_wire[8]) );
  NAND2X1 fu_ALU_fu_arch_U96 ( .A(n2201), .B(fu_ALU_fu_arch_sub_200_B_9_), .Y(
        fu_ALU_fu_arch_n260) );
  OAI211X1 fu_ALU_fu_arch_U132 ( .A0(n1778), .A1(n2093), .B0(
        fu_ALU_fu_arch_n326), .C0(fu_ALU_fu_arch_n327), .Y(fu_ALU_fu_arch_n325) );
  AOI22X1 fu_ALU_fu_arch_U57 ( .A0(n2191), .A1(fu_ALU_fu_arch_N618), .B0(n2193), .B1(fu_ALU_fu_arch_N39), .Y(fu_ALU_fu_arch_n189) );
  NAND2X1 fu_ALU_fu_arch_U69 ( .A(n1762), .B(n1754), .Y(fu_ALU_fu_arch_n210)
         );
  AOI22X1 fu_ALU_fu_arch_U310 ( .A0(n2202), .A1(fu_ALU_o1reg[8]), .B0(n2200), 
        .B1(n2168), .Y(fu_ALU_fu_arch_n552) );
  AOI221X4 U617 ( .A0(n2186), .A1(ic_socket_gcu_o1_data0_wire[5]), .B0(n2257), 
        .B1(ic_socket_ALU_o1_data0_wire[5]), .C0(n372), .Y(n368) );
  AOI22X1 fu_ALU_fu_arch_U78 ( .A0(n2191), .A1(fu_ALU_fu_arch_N616), .B0(n2193), .B1(fu_ALU_fu_arch_N37), .Y(fu_ALU_fu_arch_n223) );
  OAI22X1 fu_ALU_fu_arch_U75 ( .A0(fu_ALU_fu_arch_n208), .A1(
        fu_ALU_fu_arch_n220), .B0(fu_ALU_fu_arch_n221), .B1(n2171), .Y(
        fu_ALU_fu_arch_n219) );
  NAND2X1 fu_ALU_fu_arch_U93 ( .A(n2200), .B(fu_ALU_fu_arch_sub_200_B_4_), .Y(
        fu_ALU_fu_arch_n254) );
  OAI211X1 fu_ALU_fu_arch_U92 ( .A0(n1754), .A1(n1769), .B0(
        fu_ALU_fu_arch_n253), .C0(fu_ALU_fu_arch_n254), .Y(fu_ALU_fu_arch_n251) );
  AOI22X1 fu_ALU_fu_arch_U90 ( .A0(n2105), .A1(n1834), .B0(n2104), .B1(n1800), 
        .Y(fu_ALU_fu_arch_n246) );
  AOI22X1 fu_ALU_fu_arch_U87 ( .A0(n2191), .A1(fu_ALU_fu_arch_N615), .B0(n2193), .B1(fu_ALU_fu_arch_N36), .Y(fu_ALU_fu_arch_n239) );
  OAI22X1 fu_ALU_fu_arch_U84 ( .A0(fu_ALU_fu_arch_n234), .A1(
        fu_ALU_fu_arch_n235), .B0(fu_ALU_fu_arch_n236), .B1(n1773), .Y(
        fu_ALU_fu_arch_n233) );
  AOI22X1 fu_ALU_fu_arch_U138 ( .A0(n2191), .A1(fu_ALU_fu_arch_N614), .B0(
        n2193), .B1(fu_ALU_fu_arch_N35), .Y(fu_ALU_fu_arch_n336) );
  AOI22X1 fu_ALU_fu_arch_U127 ( .A0(n2105), .A1(n1827), .B0(n2104), .B1(n1792), 
        .Y(fu_ALU_fu_arch_n321) );
  AOI22X1 fu_ALU_fu_arch_U315 ( .A0(n2192), .A1(fu_ALU_fu_arch_N613), .B0(
        n2193), .B1(fu_ALU_fu_arch_N34), .Y(fu_ALU_fu_arch_n559) );
  OAI22X1 fu_ALU_fu_arch_U312 ( .A0(n1798), .A1(fu_ALU_fu_arch_n235), .B0(
        fu_ALU_fu_arch_n556), .B1(n1738), .Y(fu_ALU_fu_arch_n555) );
  AOI22X1 fu_ALU_fu_arch_U307 ( .A0(n2197), .A1(n2177), .B0(n2202), .B1(
        fu_ALU_fu_arch_sub_200_B_4_), .Y(fu_ALU_fu_arch_n549) );
  AOI31X1 fu_ALU_fu_arch_U306 ( .A0(fu_ALU_fu_arch_n549), .A1(
        fu_ALU_fu_arch_n550), .A2(fu_ALU_fu_arch_n551), .B0(n2106), .Y(
        fu_ALU_fu_arch_n542) );
  OAI22X1 fu_ALU_fu_arch_U303 ( .A0(fu_ALU_fu_arch_n133), .A1(
        fu_ALU_fu_arch_n544), .B0(fu_ALU_fu_arch_n137), .B1(
        fu_ALU_fu_arch_n468), .Y(fu_ALU_fu_arch_n543) );
  AOI221X4 U1158 ( .A0(n2186), .A1(ic_socket_gcu_o1_data0_wire[0]), .B0(n2257), 
        .B1(ic_socket_ALU_o1_data0_wire[0]), .C0(n613), .Y(n607) );
  OAI21X1 U1156 ( .A0(rf_BOOL_r1opcode_wire_0_), .A1(rf_BOOL_reg_0__0_), .B0(
        ic_socket_bool_o1_bus_cntrl_wire_0_), .Y(n612) );
  AOI21X1 U1155 ( .A0(rf_BOOL_r1opcode_wire_0_), .A1(n604), .B0(n612), .Y(n611) );
  AOI222X1 fu_ALU_fu_arch_U106 ( .A0(fu_ALU_fu_arch_n285), .A1(n1775), .B0(
        n1799), .B1(n2105), .C0(n1793), .C1(fu_ALU_fu_arch_n248), .Y(
        fu_ALU_fu_arch_n275) );
  AOI22X1 fu_ALU_fu_arch_U105 ( .A0(n2202), .A1(fu_ALU_o1reg[28]), .B0(n2201), 
        .B1(fu_ALU_fu_arch_sub_200_B_29_), .Y(fu_ALU_fu_arch_n282) );
  OAI21X1 fu_ALU_fu_arch_U102 ( .A0(n2172), .A1(fu_ALU_fu_arch_n275), .B0(
        fu_ALU_fu_arch_n276), .Y(fu_ALU_fu_arch_n267) );
  AOI221X2 fu_ALU_fu_arch_U101 ( .A0(n2099), .A1(n2180), .B0(
        fu_ALU_fu_arch_n175), .B1(n1739), .C0(fu_ALU_fu_arch_n274), .Y(
        fu_ALU_fu_arch_n271) );
  AOI22X1 U944 ( .A0(n2217), .A1(rf_RF_reg_3__31_), .B0(n2215), .B1(
        rf_RF_reg_1__31_), .Y(n517) );
  AOI2BB2X4 U1147 ( .B0(n604), .B1(n605), .A0N(n605), .A1N(n2111), .Y(n597) );
  AOI21X1 U1030 ( .A0(n554), .A1(inst_decoder_N121), .B0(
        inst_fetch_pc_opcode_wire_0_), .Y(n555) );
  AOI31X1 U1029 ( .A0(n1859), .A1(n536), .A2(inst_decoder_N121), .B0(n555), 
        .Y(n1134) );
  AOI21X1 U1035 ( .A0(n1859), .A1(n531), .B0(rf_BOOL_t1opcode_wire_0_), .Y(
        n560) );
  AOI31X1 U1034 ( .A0(n1859), .A1(n536), .A2(n531), .B0(n560), .Y(n1137) );
  AOI21X1 U1042 ( .A0(n1857), .A1(n553), .B0(fu_LIFTING_t1opcode_wire[0]), .Y(
        n564) );
  AOI21X1 U1040 ( .A0(n537), .A1(n1857), .B0(fu_LIFTING_t1opcode_wire[1]), .Y(
        n563) );
  AOI21X1 U1045 ( .A0(n531), .A1(n1857), .B0(fu_LIFTING_t1opcode_wire[2]), .Y(
        n565) );
  OAI21X1 U982 ( .A0(n524), .A1(n2210), .B0(n532), .Y(n1112) );
  AOI21X1 U1117 ( .A0(n1893), .A1(inst_decoder_instructionword_wire[35]), .B0(
        rf_BOOL_r1opcode_wire_0_), .Y(n589) );
  AOI31X1 U1116 ( .A0(n1893), .A1(n576), .A2(
        inst_decoder_instructionword_wire[35]), .B0(n589), .Y(n1185) );
  NAND2X1 U1059 ( .A(fu_LIFTING_in2_load_wire), .B(n2211), .Y(n569) );
  NAND2X1 U1062 ( .A(inst_fetch_ra_load_wire), .B(n2211), .Y(n570) );
  OR2X2 U1027 ( .A(n553), .B(n540), .Y(n544) );
  CLKNAND2X8 U755 ( .A(n25), .B(n2183), .Y(n250) );
  AOI211X4 U722 ( .A0(fu_LSU_t1opcode_wire[1]), .A1(n2183), .B0(n2110), .C0(
        n2247), .Y(n233) );
  AOI22X1 U315 ( .A0(n2123), .A1(rf_RF_t1data_wire[16]), .B0(
        fu_LSU_data_out[16]), .B1(n2249), .Y(n236) );
  AOI31X1 U312 ( .A0(n2185), .A1(n2111), .A2(n1826), .B0(n234), .Y(n232) );
  OAI31X4 U292 ( .A0(n220), .A1(n2183), .A2(n2110), .B0(n25), .Y(n207) );
  NAND2X1 U268 ( .A(n2123), .B(rf_RF_t1data_wire[18]), .Y(n205) );
  NAND2X1 U226 ( .A(n2123), .B(rf_RF_t1data_wire[20]), .Y(n181) );
  NAND2X1 U184 ( .A(n2123), .B(rf_RF_t1data_wire[22]), .Y(n157) );
  NAND2X1 U205 ( .A(n2123), .B(rf_RF_t1data_wire[21]), .Y(n169) );
  NAND2X1 U163 ( .A(n2123), .B(rf_RF_t1data_wire[23]), .Y(n144) );
  NAND2X1 U247 ( .A(n2123), .B(rf_RF_t1data_wire[19]), .Y(n193) );
  AOI22X1 U51 ( .A0(n2123), .A1(rf_RF_t1data_wire[28]), .B0(n29), .B1(n78), 
        .Y(n77) );
  AOI22X1 U72 ( .A0(n2123), .A1(rf_RF_t1data_wire[27]), .B0(n29), .B1(n90), 
        .Y(n89) );
  AOI22X1 U93 ( .A0(n2123), .A1(rf_RF_t1data_wire[26]), .B0(n29), .B1(n102), 
        .Y(n101) );
  OAI21X1 U453 ( .A0(n99), .A1(n250), .B0(n307), .Y(n859) );
  OAI21X1 U336 ( .A0(n24), .A1(n250), .B0(n251), .Y(n801) );
  OAI21X1 U366 ( .A0(n62), .A1(n250), .B0(n270), .Y(n814) );
  OAI21X1 U482 ( .A0(n112), .A1(n250), .B0(n318), .Y(n874) );
  OAI21X1 U424 ( .A0(n87), .A1(n250), .B0(n296), .Y(n844) );
  OAI21X1 U358 ( .A0(n35), .A1(n250), .B0(n262), .Y(n811) );
  OAI21X1 U395 ( .A0(n75), .A1(n250), .B0(n285), .Y(n829) );
  AOI21X1 U115 ( .A0(n2123), .A1(rf_RF_t1data_wire[25]), .B0(n114), .Y(n113)
         );
  AOI22X1 U137 ( .A0(n128), .A1(n129), .B0(n2123), .B1(rf_RF_t1data_wire[24]), 
        .Y(n127) );
  OAI21X1 U1149 ( .A0(n605), .A1(n2211), .B0(rf_BOOL_reg_1__0_), .Y(n606) );
  OAI21X1 U904 ( .A0(n220), .A1(n1282), .B0(n505), .Y(n1077) );
  AOI22X1 U898 ( .A0(ic_socket_gcu_o1_data0_wire[0]), .A1(n2115), .B0(
        inst_fetch_increased_pc_0_), .B1(n2116), .Y(n503) );
  OAI21X1 U897 ( .A0(n220), .A1(n264), .B0(n503), .Y(n1074) );
  AOI22X1 U1051 ( .A0(n1761), .A1(n220), .B0(n519), .B1(n2244), .Y(n1143) );
  OAI21X1 U1033 ( .A0(n559), .A1(n2211), .B0(rf_BOOL_reg_0__0_), .Y(n558) );
  OAI21X1 U1032 ( .A0(n557), .A1(n2211), .B0(n558), .Y(n1136) );
  NAND3X6 U817 ( .A(n2213), .B(n456), .C(n446), .Y(n460) );
  OAI31X4 U816 ( .A0(n470), .A1(n446), .A2(n2212), .B0(n453), .Y(n463) );
  OAI21X1 U909 ( .A0(n263), .A1(n1282), .B0(n506), .Y(n1080) );
  OAI21X1 U362 ( .A0(n263), .A1(n264), .B0(n265), .Y(n812) );
  OAI21X1 U372 ( .A0(n272), .A1(n1282), .B0(n274), .Y(n817) );
  OAI21X1 U517 ( .A0(n333), .A1(n1282), .B0(n335), .Y(n892) );
  OAI21X1 U401 ( .A0(n286), .A1(n1282), .B0(n287), .Y(n832) );
  OAI21X1 U839 ( .A0(n2213), .A1(n174), .B0(n481), .Y(n1054) );
  OAI21X1 U870 ( .A0(n2213), .A1(n491), .B0(n492), .Y(n1064) );
  OAI21X1 U833 ( .A0(n2213), .A1(n198), .B0(n479), .Y(n1052) );
  OAI21X1 U824 ( .A0(n2213), .A1(n245), .B0(n476), .Y(n1049) );
  OAI21X1 U842 ( .A0(n2213), .A1(n162), .B0(n482), .Y(n1055) );
  OAI21X1 U845 ( .A0(n2213), .A1(n150), .B0(n483), .Y(n1056) );
  OAI21X1 U836 ( .A0(n2213), .A1(n186), .B0(n480), .Y(n1053) );
  OAI21X1 U827 ( .A0(n2213), .A1(n225), .B0(n477), .Y(n1050) );
  OAI21X1 U830 ( .A0(n2213), .A1(n212), .B0(n478), .Y(n1051) );
  OAI21X1 U625 ( .A0(n375), .A1(n1282), .B0(n376), .Y(n952) );
  OAI21X1 U637 ( .A0(n375), .A1(n264), .B0(n377), .Y(n962) );
  OAI21X1 U488 ( .A0(n321), .A1(n1282), .B0(n322), .Y(n877) );
  OAI21X1 U500 ( .A0(n321), .A1(n264), .B0(n323), .Y(n887) );
  OAI21X1 U598 ( .A0(n365), .A1(n1282), .B0(n366), .Y(n937) );
  OAI21X1 U610 ( .A0(n365), .A1(n264), .B0(n367), .Y(n947) );
  OAI21X1 U430 ( .A0(n297), .A1(n1282), .B0(n298), .Y(n847) );
  OAI21X1 U544 ( .A0(n345), .A1(n1282), .B0(n346), .Y(n907) );
  OAI21X1 U556 ( .A0(n345), .A1(n264), .B0(n347), .Y(n917) );
  OAI21X1 U442 ( .A0(n297), .A1(n264), .B0(n299), .Y(n857) );
  OAI21X1 U681 ( .A0(n395), .A1(n1282), .B0(n396), .Y(n982) );
  OAI21X1 U571 ( .A0(n355), .A1(n1282), .B0(n356), .Y(n922) );
  OAI21X1 U583 ( .A0(n355), .A1(n264), .B0(n357), .Y(n932) );
  OAI21X1 U693 ( .A0(n395), .A1(n264), .B0(n397), .Y(n992) );
  OAI21X1 U459 ( .A0(n308), .A1(n1282), .B0(n309), .Y(n862) );
  OAI21X1 U471 ( .A0(n308), .A1(n264), .B0(n310), .Y(n872) );
  OAI21X1 U745 ( .A0(n2117), .A1(n1282), .B0(n410), .Y(n1028) );
  OAI21X1 U894 ( .A0(n2117), .A1(n264), .B0(n502), .Y(n1073) );
  OAI21X1 U652 ( .A0(n385), .A1(n1282), .B0(n386), .Y(n967) );
  OAI21X1 U664 ( .A0(n385), .A1(n264), .B0(n387), .Y(n977) );
  AOI21X1 U957 ( .A0(fu_LSU_t1opcode_wire[1]), .A1(n2183), .B0(n526), .Y(n528)
         );
  CLKINVX1 U1162 ( .A(inst_fetch_reset_lock), .Y(n617) );
  AOI22X1 U971 ( .A0(n498), .A1(n535), .B0(n458), .B1(n2211), .Y(n1107) );
  AOI22X1 U883 ( .A0(n498), .A1(n499), .B0(n446), .B1(n2211), .Y(n1065) );
  AOI22X1 U959 ( .A0(n498), .A1(n529), .B0(n454), .B1(n2211), .Y(n1102) );
  INVX4 fu_ALU_fu_arch_U298 ( .A(n1844), .Y(fu_ALU_fu_arch_n457) );
  AOI22X4 fu_ALU_fu_arch_U224 ( .A0(n1775), .A1(fu_ALU_fu_arch_n456), .B0(
        fu_ALU_fu_arch_n249), .B1(fu_ALU_fu_arch_n457), .Y(fu_ALU_fu_arch_n147) );
  NOR2X1 fu_ALU_fu_arch_U221 ( .A(fu_ALU_o1reg[24]), .B(n2195), .Y(
        fu_ALU_fu_arch_n455) );
  CLKNAND2X12 fu_ALU_fu_arch_U653 ( .A(n1850), .B(fu_ALU_fu_arch_n220), .Y(
        fu_ALU_fu_arch_n108) );
  AOI211X4 fu_ALU_fu_arch_U214 ( .A0(fu_ALU_fu_arch_n242), .A1(
        fu_ALU_fu_arch_n142), .B0(fu_ALU_fu_arch_n447), .C0(
        fu_ALU_fu_arch_n448), .Y(fu_ALU_fu_arch_n442) );
  AOI211X4 fu_ALU_fu_arch_U169 ( .A0(n2190), .A1(n2131), .B0(
        fu_ALU_fu_arch_n385), .C0(fu_ALU_fu_arch_n386), .Y(fu_ALU_fu_arch_n382) );
  AOI22X4 fu_ALU_fu_arch_U579 ( .A0(n2198), .A1(n2125), .B0(n1774), .B1(n2199), 
        .Y(fu_ALU_fu_arch_n592) );
  AOI22X4 fu_ALU_fu_arch_U567 ( .A0(n2198), .A1(fu_ALU_fu_arch_sub_200_B_30_), 
        .B0(n2200), .B1(fu_ALU_o1reg[31]), .Y(fu_ALU_fu_arch_n298) );
  AOI211X4 fu_ALU_fu_arch_U112 ( .A0(fu_ALU_fu_arch_sub_200_B_30_), .A1(
        fu_ALU_fu_arch_n295), .B0(fu_ALU_fu_arch_n296), .C0(
        fu_ALU_fu_arch_n297), .Y(fu_ALU_fu_arch_n294) );
  NOR2X1 fu_ALU_fu_arch_U239 ( .A(fu_ALU_o1reg[23]), .B(n2195), .Y(
        fu_ALU_fu_arch_n478) );
  AOI211X4 fu_ALU_fu_arch_U232 ( .A0(fu_ALU_fu_arch_n242), .A1(
        fu_ALU_fu_arch_n177), .B0(fu_ALU_fu_arch_n470), .C0(
        fu_ALU_fu_arch_n471), .Y(fu_ALU_fu_arch_n464) );
  OAI211X4 fu_ALU_fu_arch_U146 ( .A0(fu_ALU_fu_arch_n351), .A1(
        fu_ALU_fu_arch_n292), .B0(n2102), .C0(fu_ALU_fu_arch_n353), .Y(
        fu_ALU_fu_arch_n340) );
  OAI32X4 fu_ALU_fu_arch_U140 ( .A0(fu_ALU_fu_arch_n340), .A1(
        fu_ALU_fu_arch_n341), .A2(fu_ALU_fu_arch_n342), .B0(n1850), .B1(
        fu_ALU_fu_arch_n340), .Y(fu_ALU_fu_arch_n339) );
  AOI211X4 fu_ALU_fu_arch_U182 ( .A0(n2190), .A1(n2133), .B0(
        fu_ALU_fu_arch_n406), .C0(fu_ALU_fu_arch_n407), .Y(fu_ALU_fu_arch_n403) );
  NOR2X1 fu_ALU_fu_arch_U256 ( .A(fu_ALU_o1reg[22]), .B(n2195), .Y(
        fu_ALU_fu_arch_n497) );
  AOI211X4 fu_ALU_fu_arch_U249 ( .A0(fu_ALU_fu_arch_n242), .A1(
        fu_ALU_fu_arch_n190), .B0(fu_ALU_fu_arch_n489), .C0(
        fu_ALU_fu_arch_n490), .Y(fu_ALU_fu_arch_n484) );
  OAI211X4 fu_ALU_fu_arch_U159 ( .A0(fu_ALU_fu_arch_n372), .A1(
        fu_ALU_fu_arch_n292), .B0(n2102), .C0(fu_ALU_fu_arch_n373), .Y(
        fu_ALU_fu_arch_n361) );
  OAI32X4 fu_ALU_fu_arch_U153 ( .A0(fu_ALU_fu_arch_n361), .A1(
        fu_ALU_fu_arch_n362), .A2(fu_ALU_fu_arch_n363), .B0(n1850), .B1(
        fu_ALU_fu_arch_n361), .Y(fu_ALU_fu_arch_n360) );
  AOI211X4 fu_ALU_fu_arch_U197 ( .A0(fu_ALU_fu_arch_n242), .A1(
        fu_ALU_fu_arch_n112), .B0(fu_ALU_fu_arch_n423), .C0(
        fu_ALU_fu_arch_n424), .Y(fu_ALU_fu_arch_n418) );
  OAI22X4 fu_ALU_fu_arch_U279 ( .A0(fu_ALU_fu_arch_n135), .A1(n2106), .B0(
        fu_ALU_fu_arch_n519), .B1(n2203), .Y(fu_ALU_fu_arch_n511) );
  AOI211X4 fu_ALU_fu_arch_U266 ( .A0(fu_ALU_fu_arch_n333), .A1(n1882), .B0(
        fu_ALU_fu_arch_n508), .C0(fu_ALU_fu_arch_n509), .Y(fu_ALU_fu_arch_n503) );
  NOR2X1 fu_ALU_fu_arch_U265 ( .A(n2143), .B(n2195), .Y(fu_ALU_fu_arch_n507)
         );
  NAND4X4 fu_ALU_fu_arch_U689 ( .A(fu_ALU_fu_arch_n446), .B(
        fu_ALU_fu_arch_n767), .C(fu_ALU_fu_arch_n412), .D(fu_ALU_fu_arch_n487), 
        .Y(fu_ALU_fu_arch_n534) );
  AOI211X4 fu_ALU_fu_arch_U284 ( .A0(fu_ALU_fu_arch_n242), .A1(
        fu_ALU_fu_arch_n214), .B0(fu_ALU_fu_arch_n525), .C0(
        fu_ALU_fu_arch_n526), .Y(fu_ALU_fu_arch_n520) );
  AOI211X4 fu_ALU_fu_arch_U322 ( .A0(fu_ALU_fu_arch_n240), .A1(
        fu_ALU_fu_arch_n229), .B0(fu_ALU_fu_arch_n567), .C0(
        fu_ALU_fu_arch_n568), .Y(fu_ALU_fu_arch_n560) );
  NOR2X1 fu_ALU_fu_arch_U320 ( .A(n2147), .B(n2195), .Y(fu_ALU_fu_arch_n566)
         );
  AOI21X4 fu_ALU_fu_arch_U351 ( .A0(n2105), .A1(fu_ALU_fu_arch_n592), .B0(
        fu_ALU_fu_arch_n591), .Y(fu_ALU_fu_arch_n316) );
  AOI211X4 fu_ALU_fu_arch_U341 ( .A0(fu_ALU_fu_arch_n240), .A1(
        fu_ALU_fu_arch_n328), .B0(fu_ALU_fu_arch_n584), .C0(
        fu_ALU_fu_arch_n585), .Y(fu_ALU_fu_arch_n577) );
  NOR2X1 fu_ALU_fu_arch_U340 ( .A(n2149), .B(n2195), .Y(fu_ALU_fu_arch_n583)
         );
  OAI211X2 fu_ALU_fu_arch_U456 ( .A0(fu_ALU_fu_arch_n522), .A1(n2199), .B0(
        fu_ALU_fu_arch_n517), .C0(fu_ALU_fu_arch_n572), .Y(fu_ALU_fu_arch_n669) );
  OAI222X4 fu_ALU_fu_arch_U373 ( .A0(n2106), .A1(fu_ALU_fu_arch_n131), .B0(
        fu_ALU_fu_arch_n468), .B1(fu_ALU_fu_arch_n519), .C0(n2203), .C1(
        fu_ALU_fu_arch_n135), .Y(fu_ALU_fu_arch_n606) );
  AOI211X4 fu_ALU_fu_arch_U359 ( .A0(fu_ALU_fu_arch_n240), .A1(
        fu_ALU_fu_arch_n539), .B0(fu_ALU_fu_arch_n599), .C0(
        fu_ALU_fu_arch_n600), .Y(fu_ALU_fu_arch_n594) );
  NOR2X1 fu_ALU_fu_arch_U391 ( .A(n2152), .B(n2195), .Y(fu_ALU_fu_arch_n620)
         );
  AOI211X4 fu_ALU_fu_arch_U382 ( .A0(fu_ALU_fu_arch_n333), .A1(n1840), .B0(
        fu_ALU_fu_arch_n613), .C0(fu_ALU_fu_arch_n614), .Y(fu_ALU_fu_arch_n609) );
  OAI2B11X2 fu_ALU_fu_arch_U397 ( .A1N(n2153), .A0(fu_ALU_fu_arch_n629), .B0(
        fu_ALU_fu_arch_n630), .C0(n2102), .Y(fu_ALU_fu_arch_n628) );
  AOI211X4 fu_ALU_fu_arch_U396 ( .A0(fu_ALU_fu_arch_n612), .A1(
        fu_ALU_fu_arch_n277), .B0(fu_ALU_fu_arch_n627), .C0(
        fu_ALU_fu_arch_n628), .Y(fu_ALU_fu_arch_n625) );
  AOI211X4 fu_ALU_fu_arch_U414 ( .A0(fu_ALU_fu_arch_n612), .A1(
        fu_ALU_fu_arch_n304), .B0(fu_ALU_fu_arch_n643), .C0(
        fu_ALU_fu_arch_n644), .Y(fu_ALU_fu_arch_n641) );
  AOI21X6 fu_ALU_fu_arch_U468 ( .A0(n2200), .A1(fu_ALU_fu_arch_sub_200_B_14_), 
        .B0(fu_ALU_fu_arch_n673), .Y(fu_ALU_fu_arch_n133) );
  NOR2X1 fu_ALU_fu_arch_U467 ( .A(n2156), .B(n2195), .Y(fu_ALU_fu_arch_n672)
         );
  NOR4X4 fu_ALU_fu_arch_U12 ( .A(fu_ALU_fu_arch_n113), .B(fu_ALU_fu_arch_n114), 
        .C(fu_ALU_fu_arch_n115), .D(fu_ALU_fu_arch_n116), .Y(
        fu_ALU_fu_arch_n109) );
  NOR4X4 fu_ALU_fu_arch_U31 ( .A(fu_ALU_fu_arch_n143), .B(fu_ALU_fu_arch_n144), 
        .C(fu_ALU_fu_arch_n145), .D(fu_ALU_fu_arch_n146), .Y(
        fu_ALU_fu_arch_n140) );
  AOI221X2 fu_ALU_fu_arch_U43 ( .A0(n1892), .A1(n1834), .B0(n1854), .B1(n1800), 
        .C0(fu_ALU_fu_arch_n165), .Y(fu_ALU_fu_arch_n160) );
  NOR4X4 fu_ALU_fu_arch_U64 ( .A(fu_ALU_fu_arch_n200), .B(fu_ALU_fu_arch_n201), 
        .C(fu_ALU_fu_arch_n202), .D(fu_ALU_fu_arch_n203), .Y(
        fu_ALU_fu_arch_n196) );
  OAI211X4 fu_ALU_fu_arch_U639 ( .A0(n2171), .A1(n2199), .B0(
        fu_ALU_fu_arch_n758), .C0(fu_ALU_fu_arch_n689), .Y(fu_ALU_fu_arch_n217) );
  AOI32X1 fu_ALU_fu_arch_U91 ( .A0(fu_ALU_fu_arch_n249), .A1(n2197), .A2(
        fu_ALU_o1reg[3]), .B0(fu_ALU_fu_arch_n251), .B1(fu_ALU_fu_arch_n249), 
        .Y(fu_ALU_fu_arch_n245) );
  OAI31X4 fu_ALU_fu_arch_U602 ( .A0(fu_ALU_fu_arch_n737), .A1(
        fu_ALU_fu_arch_n607), .A2(fu_ALU_fu_arch_n220), .B0(
        fu_ALU_fu_arch_n738), .Y(ic_socket_ALU_o1_data0_wire[0]) );
  NOR3X2 fu_ALU_fu_arch_U108 ( .A(n2124), .B(n2195), .C(n1739), .Y(
        fu_ALU_fu_arch_n289) );
  AOI22X1 U1098 ( .A0(n2207), .A1(n578), .B0(n67), .B1(n2206), .Y(n1177) );
  AOI22X1 U1100 ( .A0(n2207), .A1(n579), .B0(n513), .B1(n2206), .Y(n1178) );
  OAI2B2X1 U1031 ( .A1N(inst_fetch_pc_load_wire), .A0(n2210), .B0(n556), .B1(
        n531), .Y(n1135) );
  MX2X1 U1078 ( .A(inst_decoder_instructionword_wire[16]), .B(
        ic_simm_B1_wire[10]), .S0(n2206), .Y(n1157) );
  MX2X1 U1089 ( .A(inst_decoder_instructionword_wire[17]), .B(
        ic_simm_B1_wire[11]), .S0(n2206), .Y(n1168) );
  MX2X1 U1079 ( .A(inst_decoder_instructionword_wire[14]), .B(
        ic_simm_B1_wire[8]), .S0(n2206), .Y(n1158) );
  MX2X1 U1088 ( .A(inst_decoder_instructionword_wire[15]), .B(
        ic_simm_B1_wire[9]), .S0(n2206), .Y(n1167) );
  MX2X1 U1087 ( .A(inst_decoder_instructionword_wire[13]), .B(
        ic_simm_B1_wire[7]), .S0(n2206), .Y(n1166) );
  MX2X1 U1071 ( .A(inst_decoder_instructionword_wire[30]), .B(
        ic_simm_B1_wire[24]), .S0(n2206), .Y(n1150) );
  MX2X1 U1069 ( .A(inst_decoder_instructionword_wire[34]), .B(
        ic_simm_B1_wire[28]), .S0(n2206), .Y(n1148) );
  MX2X1 U1076 ( .A(inst_decoder_instructionword_wire[20]), .B(
        ic_simm_B1_wire[14]), .S0(n2206), .Y(n1155) );
  MX2X1 U1077 ( .A(inst_decoder_instructionword_wire[18]), .B(
        ic_simm_B1_wire[12]), .S0(n2206), .Y(n1156) );
  MX2X1 U1090 ( .A(inst_decoder_instructionword_wire[19]), .B(
        ic_simm_B1_wire[13]), .S0(n2206), .Y(n1169) );
  MX2X1 U1075 ( .A(inst_decoder_instructionword_wire[22]), .B(
        ic_simm_B1_wire[16]), .S0(n2206), .Y(n1154) );
  MX2X1 U1091 ( .A(inst_decoder_instructionword_wire[21]), .B(
        ic_simm_B1_wire[15]), .S0(n2206), .Y(n1170) );
  MX2X1 U1095 ( .A(inst_decoder_instructionword_wire[29]), .B(
        ic_simm_B1_wire[23]), .S0(n2206), .Y(n1174) );
  MX2X1 U1093 ( .A(inst_decoder_instructionword_wire[25]), .B(
        ic_simm_B1_wire[19]), .S0(n2206), .Y(n1172) );
  MX2X1 U1096 ( .A(inst_decoder_instructionword_wire[31]), .B(
        ic_simm_B1_wire[25]), .S0(n2206), .Y(n1175) );
  MX2X1 U1074 ( .A(inst_decoder_instructionword_wire[24]), .B(
        ic_simm_B1_wire[18]), .S0(n2206), .Y(n1153) );
  MX2X1 U1080 ( .A(inst_decoder_instructionword_wire[12]), .B(
        ic_simm_B1_wire[6]), .S0(n2206), .Y(n1159) );
  MX2X1 U1086 ( .A(inst_decoder_instructionword_wire[11]), .B(
        ic_simm_B1_wire[5]), .S0(n2206), .Y(n1165) );
  MX2X1 U1073 ( .A(inst_decoder_instructionword_wire[26]), .B(
        ic_simm_B1_wire[20]), .S0(n2206), .Y(n1152) );
  MX2X1 U1097 ( .A(inst_decoder_instructionword_wire[33]), .B(
        ic_simm_B1_wire[27]), .S0(n2206), .Y(n1176) );
  MX2X1 U1092 ( .A(inst_decoder_instructionword_wire[23]), .B(
        ic_simm_B1_wire[17]), .S0(n2206), .Y(n1171) );
  MX2X1 U1085 ( .A(inst_decoder_instructionword_wire[9]), .B(
        ic_simm_B1_wire[3]), .S0(n2206), .Y(n1164) );
  MX2X1 U1081 ( .A(inst_decoder_instructionword_wire[10]), .B(
        ic_simm_B1_wire[4]), .S0(n2206), .Y(n1160) );
  MX2X1 U1072 ( .A(inst_decoder_instructionword_wire[28]), .B(
        ic_simm_B1_wire[22]), .S0(n2206), .Y(n1151) );
  MX2X1 U1094 ( .A(inst_decoder_instructionword_wire[27]), .B(
        ic_simm_B1_wire[21]), .S0(n2206), .Y(n1173) );
  OAI22X1 U1036 ( .A0(inst_decoder_N121), .A1(n556), .B0(n2210), .B1(n561), 
        .Y(n1138) );
  OAI21X1 U1103 ( .A0(n2210), .A1(n1750), .B0(n2206), .Y(n1179) );
  AOI31X1 U1041 ( .A0(n1857), .A1(n536), .A2(n553), .B0(n564), .Y(n1140) );
  AOI21X1 U1039 ( .A0(n1857), .A1(n531), .B0(n563), .Y(n1139) );
  AOI21X1 U1044 ( .A0(n1857), .A1(n537), .B0(n565), .Y(n1141) );
  OAI21X1 U1113 ( .A0(n2210), .A1(n1748), .B0(n583), .Y(n1183) );
  OAI22X1 U1015 ( .A0(n549), .A1(n548), .B0(n538), .B1(n542), .Y(n1130) );
  OAI22X1 U1055 ( .A0(n2210), .A1(n521), .B0(n567), .B1(n568), .Y(n1144) );
  MX2X1 U1070 ( .A(inst_decoder_instructionword_wire[32]), .B(
        ic_simm_B1_wire[26]), .S0(n574), .Y(n1149) );
  OAI2B2X1 U1115 ( .A1N(n2186), .A0(n2210), .B0(
        inst_decoder_instructionword_wire[35]), .B1(n588), .Y(n1184) );
  AOI22X4 U649 ( .A0(n2185), .A1(n1808), .B0(fu_LSU_o1shadow_reg_3_), .B1(n132), .Y(n191) );
  AOI22X4 U568 ( .A0(n2185), .A1(n1818), .B0(fu_LSU_o1shadow_reg_6_), .B1(n132), .Y(n155) );
  AOI22X4 U541 ( .A0(n2185), .A1(n1814), .B0(fu_LSU_o1shadow_reg_7_), .B1(n132), .Y(n141) );
  AOI22X4 U595 ( .A0(n2185), .A1(n1821), .B0(fu_LSU_o1shadow_reg_5_), .B1(n132), .Y(n167) );
  AOI22X4 U622 ( .A0(n2185), .A1(n1825), .B0(fu_LSU_o1shadow_reg_4_), .B1(n132), .Y(n179) );
  AOI22X4 U678 ( .A0(fu_LSU_o1load_wire), .A1(n1810), .B0(
        fu_LSU_o1shadow_reg_2_), .B1(n132), .Y(n203) );
  MX2X1 U32 ( .A(n1861), .B(n2128), .S0(n2252), .Y(n662) );
  MX2X1 U11 ( .A(n1862), .B(n2126), .S0(n2252), .Y(n652) );
  MX2X1 U930 ( .A(n1860), .B(n2180), .S0(n2252), .Y(n1090) );
  MX2X1 U53 ( .A(rf_RF_t1data_wire[28]), .B(n2130), .S0(n2253), .Y(n672) );
  MX2X1 U74 ( .A(rf_RF_t1data_wire[27]), .B(n2131), .S0(n2252), .Y(n682) );
  MX2X1 U96 ( .A(rf_RF_t1data_wire[26]), .B(n2133), .S0(n2253), .Y(n692) );
  MX2X1 U118 ( .A(rf_RF_t1data_wire[25]), .B(n2135), .S0(n2253), .Y(n702) );
  MX2X1 U142 ( .A(rf_RF_t1data_wire[24]), .B(n2137), .S0(n2252), .Y(n712) );
  MX2X1 U165 ( .A(rf_RF_t1data_wire[23]), .B(n2139), .S0(n2252), .Y(n722) );
  AOI22X1 U961 ( .A0(n500), .A1(n220), .B0(n529), .B1(n501), .Y(n1103) );
  AOI2BB2X1 U1008 ( .B0(n2225), .B1(n220), .A0N(rf_RF_reg_4__0_), .A1N(n2226), 
        .Y(n1127) );
  MX2X1 U186 ( .A(rf_RF_t1data_wire[22]), .B(n2141), .S0(n2253), .Y(n732) );
  MX2X1 U207 ( .A(rf_RF_t1data_wire[21]), .B(n2143), .S0(n2253), .Y(n742) );
  OAI21X1 U947 ( .A0(n519), .A1(n2255), .B0(n520), .Y(n1098) );
  MX2X1 U228 ( .A(rf_RF_t1data_wire[20]), .B(n2145), .S0(n2252), .Y(n752) );
  MX2X1 U994 ( .A(n1779), .B(n2111), .S0(n2098), .Y(n1121) );
  MX2X1 U249 ( .A(rf_RF_t1data_wire[19]), .B(n2147), .S0(n2252), .Y(n762) );
  MX2X1 U271 ( .A(rf_RF_t1data_wire[18]), .B(n2149), .S0(n2253), .Y(n772) );
  OAI21X1 U529 ( .A0(n333), .A1(n264), .B0(n336), .Y(n902) );
  AOI21X1 U861 ( .A0(ic_socket_lsu_o1_data0_wire[28]), .A1(n2212), .B0(n2119), 
        .Y(n488) );
  OAI21X1 U860 ( .A0(n453), .A1(n437), .B0(n488), .Y(n1061) );
  AOI21X1 U849 ( .A0(ic_socket_lsu_o1_data0_wire[24]), .A1(n2212), .B0(n2119), 
        .Y(n484) );
  OAI21X1 U848 ( .A0(n453), .A1(n421), .B0(n484), .Y(n1057) );
  AOI21X1 U864 ( .A0(ic_socket_lsu_o1_data0_wire[29]), .A1(n2212), .B0(n2119), 
        .Y(n489) );
  OAI21X1 U863 ( .A0(n453), .A1(n440), .B0(n489), .Y(n1062) );
  AOI21X1 U852 ( .A0(ic_socket_lsu_o1_data0_wire[25]), .A1(n2212), .B0(n2119), 
        .Y(n485) );
  OAI21X1 U851 ( .A0(n453), .A1(n428), .B0(n485), .Y(n1058) );
  AOI21X1 U858 ( .A0(ic_socket_lsu_o1_data0_wire[27]), .A1(n2212), .B0(n2119), 
        .Y(n487) );
  OAI21X1 U857 ( .A0(n453), .A1(n434), .B0(n487), .Y(n1060) );
  AOI21X1 U867 ( .A0(ic_socket_lsu_o1_data0_wire[30]), .A1(n2212), .B0(n2119), 
        .Y(n490) );
  OAI21X1 U866 ( .A0(n453), .A1(n443), .B0(n490), .Y(n1063) );
  AOI21X1 U855 ( .A0(ic_socket_lsu_o1_data0_wire[26]), .A1(n2212), .B0(n2119), 
        .Y(n486) );
  OAI21X1 U854 ( .A0(n453), .A1(n431), .B0(n486), .Y(n1059) );
  MX2X1 U293 ( .A(rf_RF_t1data_wire[17]), .B(n2150), .S0(n2253), .Y(n782) );
  AOI21X1 U840 ( .A0(n2118), .A1(fu_LSU_data_in[21]), .B0(n2119), .Y(n481) );
  AOI21X1 U871 ( .A0(n2118), .A1(fu_LSU_data_in[31]), .B0(n2119), .Y(n492) );
  AOI21X1 U834 ( .A0(n2118), .A1(fu_LSU_data_in[19]), .B0(n2119), .Y(n479) );
  AOI21X1 U825 ( .A0(n2118), .A1(fu_LSU_data_in[16]), .B0(n2119), .Y(n476) );
  AOI21X1 U843 ( .A0(n2118), .A1(fu_LSU_data_in[22]), .B0(n2119), .Y(n482) );
  AOI21X1 U846 ( .A0(n2118), .A1(fu_LSU_data_in[23]), .B0(n2119), .Y(n483) );
  AOI21X1 U837 ( .A0(n2118), .A1(fu_LSU_data_in[20]), .B0(n2119), .Y(n480) );
  AOI21X1 U828 ( .A0(n2118), .A1(fu_LSU_data_in[17]), .B0(n2119), .Y(n477) );
  AOI21X1 U831 ( .A0(n2118), .A1(fu_LSU_data_in[18]), .B0(n2119), .Y(n478) );
  MX2X1 U915 ( .A(fu_LSU_addr[12]), .B(rf_RF_t1data_wire[14]), .S0(n2113), .Y(
        n1083) );
  MX2X1 U913 ( .A(rf_RF_t1data_wire[14]), .B(n2179), .S0(n2252), .Y(n1081) );
  OAI21X1 U702 ( .A0(n2255), .A1(n403), .B0(n404), .Y(n993) );
  MX2X1 U767 ( .A(n2110), .B(fu_ALU_fu_arch_sub_200_A_1_), .S0(n2253), .Y(
        n1031) );
  MX2X1 U318 ( .A(rf_RF_t1data_wire[16]), .B(n2152), .S0(n2252), .Y(n792) );
  MX2X1 U376 ( .A(fu_LSU_addr[11]), .B(n1823), .S0(n2113), .Y(n820) );
  MX2X1 U374 ( .A(n1823), .B(n2156), .S0(n2252), .Y(n818) );
  OAI21X1 U619 ( .A0(n2254), .A1(n373), .B0(n374), .Y(n948) );
  OAI21X1 U480 ( .A0(n2255), .A1(n316), .B0(n317), .Y(n873) );
  OAI21X1 U592 ( .A0(n2255), .A1(n363), .B0(n364), .Y(n933) );
  MX2X1 U405 ( .A(fu_LSU_addr[10]), .B(n1820), .S0(n2113), .Y(n835) );
  MX2X1 U403 ( .A(n1820), .B(n2158), .S0(n2253), .Y(n833) );
  OAI21X1 U565 ( .A0(n2255), .A1(n353), .B0(n354), .Y(n918) );
  MX2X1 U629 ( .A(fu_LSU_addr[2]), .B(n1825), .S0(n2113), .Y(n955) );
  MX2X1 U340 ( .A(rf_RF_t1data_wire[15]), .B(n2154), .S0(n2252), .Y(n802) );
  MX2X1 U492 ( .A(fu_LSU_addr[7]), .B(n1812), .S0(n2113), .Y(n880) );
  OAI21X1 U509 ( .A0(n2255), .A1(n329), .B0(n330), .Y(n888) );
  MX2X1 U602 ( .A(fu_LSU_addr[3]), .B(n1821), .S0(n2113), .Y(n940) );
  MX2X1 U490 ( .A(n1812), .B(n2163), .S0(n2252), .Y(n878) );
  OAI21X1 U538 ( .A0(n2255), .A1(n342), .B0(n343), .Y(n903) );
  OAI21X1 U673 ( .A0(n2254), .A1(n393), .B0(n394), .Y(n978) );
  MX2X1 U521 ( .A(fu_LSU_addr[6]), .B(rf_RF_t1data_wire[8]), .S0(n2113), .Y(
        n895) );
  MX2X1 U548 ( .A(fu_LSU_addr[5]), .B(n1814), .S0(n2113), .Y(n910) );
  MX2X1 U519 ( .A(rf_RF_t1data_wire[8]), .B(n2165), .S0(n2253), .Y(n893) );
  MX2X1 U546 ( .A(n1814), .B(n2167), .S0(n2252), .Y(n908) );
  MX2X1 U575 ( .A(fu_LSU_addr[4]), .B(n1818), .S0(n2113), .Y(n925) );
  MX2X1 U573 ( .A(n1818), .B(n2169), .S0(n2253), .Y(n923) );
  OAI21X1 U451 ( .A0(n2255), .A1(n305), .B0(n306), .Y(n858) );
  MX2X1 U434 ( .A(fu_LSU_addr[9]), .B(rf_RF_t1data_wire[11]), .S0(n2113), .Y(
        n850) );
  MX2X1 U432 ( .A(rf_RF_t1data_wire[11]), .B(n2160), .S0(n2252), .Y(n848) );
  MX2X1 U685 ( .A(fu_LSU_addr[0]), .B(n1810), .S0(n2113), .Y(n985) );
  MX2X1 U683 ( .A(n1810), .B(n2176), .S0(n2252), .Y(n983) );
  OAI21X1 U646 ( .A0(n2254), .A1(n383), .B0(n384), .Y(n963) );
  MX2X1 U656 ( .A(fu_LSU_addr[1]), .B(n1808), .S0(n2113), .Y(n970) );
  MX2X1 U463 ( .A(fu_LSU_addr[8]), .B(n1816), .S0(n2113), .Y(n865) );
  MX2X1 U461 ( .A(n1816), .B(n2162), .S0(n2253), .Y(n863) );
  MX2X1 U1237 ( .A(inst_fetch_N59), .B(inst_fetch_reset_cntr_13_), .S0(n2205), 
        .Y(n1255) );
  MX2X1 U1222 ( .A(inst_fetch_N62), .B(inst_fetch_reset_cntr_16_), .S0(n2204), 
        .Y(n1240) );
  MX2X1 U1224 ( .A(inst_fetch_N58), .B(inst_fetch_reset_cntr_12_), .S0(n2204), 
        .Y(n1242) );
  MX2X1 U1231 ( .A(inst_fetch_N47), .B(inst_fetch_reset_cntr_1_), .S0(n2205), 
        .Y(n1249) );
  MX2X1 U1242 ( .A(inst_fetch_N69), .B(inst_fetch_reset_cntr_23_), .S0(n2205), 
        .Y(n1260) );
  MX2X1 U1233 ( .A(inst_fetch_N51), .B(inst_fetch_reset_cntr_5_), .S0(n2205), 
        .Y(n1251) );
  MX2X1 U1239 ( .A(inst_fetch_N63), .B(inst_fetch_reset_cntr_17_), .S0(n2205), 
        .Y(n1257) );
  MX2X1 U1218 ( .A(inst_fetch_N70), .B(inst_fetch_reset_cntr_24_), .S0(n2204), 
        .Y(n1236) );
  MX2X1 U1227 ( .A(inst_fetch_N52), .B(inst_fetch_reset_cntr_6_), .S0(n2204), 
        .Y(n1245) );
  MX2X1 U1234 ( .A(inst_fetch_N53), .B(inst_fetch_reset_cntr_7_), .S0(n2205), 
        .Y(n1252) );
  MX2X1 U1219 ( .A(inst_fetch_N68), .B(inst_fetch_reset_cntr_22_), .S0(n2204), 
        .Y(n1237) );
  MX2X1 U1235 ( .A(inst_fetch_N55), .B(inst_fetch_reset_cntr_9_), .S0(n2205), 
        .Y(n1253) );
  MX2X1 U1232 ( .A(inst_fetch_N49), .B(inst_fetch_reset_cntr_3_), .S0(n2205), 
        .Y(n1250) );
  MX2X1 U1220 ( .A(inst_fetch_N66), .B(inst_fetch_reset_cntr_20_), .S0(n2204), 
        .Y(n1238) );
  MX2X1 U1229 ( .A(inst_fetch_N48), .B(inst_fetch_reset_cntr_2_), .S0(n2205), 
        .Y(n1247) );
  MX2X1 U1238 ( .A(inst_fetch_N61), .B(inst_fetch_reset_cntr_15_), .S0(n2205), 
        .Y(n1256) );
  MX2X1 U1240 ( .A(inst_fetch_N65), .B(inst_fetch_reset_cntr_19_), .S0(n2205), 
        .Y(n1258) );
  MX2X1 U1241 ( .A(inst_fetch_N67), .B(inst_fetch_reset_cntr_21_), .S0(n2205), 
        .Y(n1259) );
  MX2X1 U1221 ( .A(inst_fetch_N64), .B(inst_fetch_reset_cntr_18_), .S0(n2204), 
        .Y(n1239) );
  MX2X1 U1223 ( .A(inst_fetch_N60), .B(inst_fetch_reset_cntr_14_), .S0(n2204), 
        .Y(n1241) );
  MX2X1 U1226 ( .A(inst_fetch_N54), .B(inst_fetch_reset_cntr_8_), .S0(n2204), 
        .Y(n1244) );
  MX2X1 U1228 ( .A(inst_fetch_N50), .B(inst_fetch_reset_cntr_4_), .S0(n2204), 
        .Y(n1246) );
  MX2X1 U1225 ( .A(inst_fetch_N56), .B(inst_fetch_reset_cntr_10_), .S0(n2204), 
        .Y(n1243) );
  MX2X1 U1236 ( .A(inst_fetch_N57), .B(inst_fetch_reset_cntr_11_), .S0(n2205), 
        .Y(n1254) );
  OAI22X1 U969 ( .A0(n2210), .A1(n533), .B0(n534), .B1(n1751), .Y(n1106) );
  OAI22X1 U973 ( .A0(n2183), .A1(n534), .B0(n2210), .B1(n535), .Y(n1108) );
  OAI221X1 U956 ( .A0(n526), .A1(n527), .B0(n528), .B1(fu_LSU_t1opcode_wire[2]), .C0(n2113), .Y(n525) );
  OAI2BB1X1 U955 ( .A0N(fu_LSU_status_addr_reg_0__2_), .A1N(n2211), .B0(n525), 
        .Y(n1101) );
  AOI31X1 U1161 ( .A0(n614), .A1(n615), .A2(n616), .B0(n617), .Y(n1191) );
  MX2X1 U992 ( .A(fu_ALU_t1opcode_wire[3]), .B(fu_ALU_opc1reg[3]), .S0(n2252), 
        .Y(n1119) );
  MX2X1 U988 ( .A(fu_ALU_t1opcode_wire[0]), .B(fu_ALU_opc1reg[0]), .S0(n2252), 
        .Y(n1115) );
  MX2X1 U990 ( .A(fu_ALU_t1opcode_wire[1]), .B(fu_ALU_opc1reg[1]), .S0(n2252), 
        .Y(n1117) );
  MX2X1 U986 ( .A(fu_ALU_t1opcode_wire[2]), .B(fu_ALU_opc1reg[2]), .S0(n2252), 
        .Y(n1113) );
  OAI2B2X1 U981 ( .A1N(fu_LSU_mem_en_x[0]), .A0(n2210), .B0(n2211), .B1(
        fu_LSU_t1load_wire), .Y(n1111) );
  AOI2BB2X1 U953 ( .B0(n459), .B1(n2211), .A0N(n2211), .A1N(
        fu_LSU_status_addr_reg_0__2_), .Y(n1100) );
  AOI2BB2X1 U968 ( .B0(n2210), .B1(n533), .A0N(fu_LSU_status_addr_reg_1__4_), 
        .A1N(n2210), .Y(n1105) );
  MX2X1 U1214 ( .A(inst_decoder_N121), .B(imem_data[1]), .S0(n2208), .Y(n1232)
         );
  MX2X1 U1175 ( .A(inst_decoder_instructionword_wire[40]), .B(imem_data[40]), 
        .S0(n2209), .Y(n1193) );
  MX2X1 U1200 ( .A(inst_decoder_instructionword_wire[15]), .B(imem_data[15]), 
        .S0(n2209), .Y(n1218) );
  MX2X1 U1181 ( .A(inst_decoder_instructionword_wire[34]), .B(imem_data[34]), 
        .S0(n2209), .Y(n1199) );
  MX2X1 U1183 ( .A(inst_decoder_instructionword_wire[32]), .B(imem_data[32]), 
        .S0(n2209), .Y(n1201) );
  MX2X1 U1185 ( .A(inst_decoder_instructionword_wire[30]), .B(imem_data[30]), 
        .S0(n2209), .Y(n1203) );
  MX2X1 U1196 ( .A(inst_decoder_instructionword_wire[19]), .B(imem_data[19]), 
        .S0(n2209), .Y(n1214) );
  MX2X1 U1176 ( .A(inst_decoder_instructionword_wire[39]), .B(imem_data[39]), 
        .S0(n2209), .Y(n1194) );
  MX2X1 U1191 ( .A(inst_decoder_instructionword_wire[24]), .B(imem_data[24]), 
        .S0(n2209), .Y(n1209) );
  MX2X1 U1199 ( .A(inst_decoder_instructionword_wire[16]), .B(imem_data[16]), 
        .S0(n2209), .Y(n1217) );
  MX2X1 U1198 ( .A(inst_decoder_instructionword_wire[17]), .B(imem_data[17]), 
        .S0(n2209), .Y(n1216) );
  MX2X1 U1187 ( .A(inst_decoder_instructionword_wire[28]), .B(imem_data[28]), 
        .S0(n2209), .Y(n1205) );
  MX2X1 U1205 ( .A(inst_decoder_instructionword_wire[10]), .B(imem_data[10]), 
        .S0(n2209), .Y(n1223) );
  MX2X1 U1204 ( .A(inst_decoder_instructionword_wire[11]), .B(imem_data[11]), 
        .S0(n2209), .Y(n1222) );
  MX2X1 U1203 ( .A(inst_decoder_instructionword_wire[12]), .B(imem_data[12]), 
        .S0(n2209), .Y(n1221) );
  MX2X1 U1202 ( .A(inst_decoder_instructionword_wire[13]), .B(imem_data[13]), 
        .S0(n2209), .Y(n1220) );
  MX2X1 U1201 ( .A(inst_decoder_instructionword_wire[14]), .B(imem_data[14]), 
        .S0(n2209), .Y(n1219) );
  MX2X1 U1194 ( .A(inst_decoder_instructionword_wire[21]), .B(imem_data[21]), 
        .S0(n2209), .Y(n1212) );
  MX2X1 U1193 ( .A(inst_decoder_instructionword_wire[22]), .B(imem_data[22]), 
        .S0(n2209), .Y(n1211) );
  MX2X1 U1188 ( .A(inst_decoder_instructionword_wire[27]), .B(imem_data[27]), 
        .S0(n2209), .Y(n1206) );
  MX2X1 U1197 ( .A(inst_decoder_instructionword_wire[18]), .B(imem_data[18]), 
        .S0(n2209), .Y(n1215) );
  MX2X1 U1189 ( .A(inst_decoder_instructionword_wire[26]), .B(imem_data[26]), 
        .S0(n2209), .Y(n1207) );
  MX2X1 U1195 ( .A(inst_decoder_instructionword_wire[20]), .B(imem_data[20]), 
        .S0(n2209), .Y(n1213) );
  MX2X1 U1192 ( .A(inst_decoder_instructionword_wire[23]), .B(imem_data[23]), 
        .S0(n2209), .Y(n1210) );
  MX2X1 U1180 ( .A(inst_decoder_instructionword_wire[35]), .B(imem_data[35]), 
        .S0(n2208), .Y(n1198) );
  MX2X1 U1213 ( .A(inst_decoder_N230), .B(imem_data[2]), .S0(n2208), .Y(n1231)
         );
  MX2X1 U1211 ( .A(inst_decoder_instructionword_wire[4]), .B(imem_data[4]), 
        .S0(n2208), .Y(n1229) );
  MX2X1 U1179 ( .A(inst_decoder_instructionword_wire[36]), .B(imem_data[36]), 
        .S0(n2208), .Y(n1197) );
  MX2X1 U1212 ( .A(inst_decoder_N232), .B(imem_data[3]), .S0(n2208), .Y(n1230)
         );
  MX2X1 U1182 ( .A(inst_decoder_instructionword_wire[33]), .B(imem_data[33]), 
        .S0(n2208), .Y(n1200) );
  MX2X1 U1184 ( .A(inst_decoder_instructionword_wire[31]), .B(imem_data[31]), 
        .S0(n2208), .Y(n1202) );
  MX2X1 U1215 ( .A(inst_decoder_N119), .B(imem_data[0]), .S0(n2208), .Y(n1233)
         );
  MX2X1 U1178 ( .A(inst_decoder_instructionword_wire[37]), .B(imem_data[37]), 
        .S0(n2208), .Y(n1196) );
  MX2X1 U1207 ( .A(inst_decoder_instructionword_wire[8]), .B(imem_data[8]), 
        .S0(n2208), .Y(n1225) );
  MX2X1 U1190 ( .A(inst_decoder_instructionword_wire[25]), .B(imem_data[25]), 
        .S0(n2208), .Y(n1208) );
  MX2X1 U1186 ( .A(inst_decoder_instructionword_wire[29]), .B(imem_data[29]), 
        .S0(n2208), .Y(n1204) );
  MX2X1 U1174 ( .A(inst_decoder_instructionword_wire[41]), .B(imem_data[41]), 
        .S0(n2208), .Y(n1192) );
  MX2X1 U1208 ( .A(inst_decoder_instructionword_wire[7]), .B(imem_data[7]), 
        .S0(n2208), .Y(n1226) );
  MX2X1 U1177 ( .A(inst_decoder_instructionword_wire[38]), .B(imem_data[38]), 
        .S0(n2208), .Y(n1195) );
  MX2X1 U1206 ( .A(inst_decoder_instructionword_wire[9]), .B(imem_data[9]), 
        .S0(n2208), .Y(n1224) );
  MX2X1 U1210 ( .A(inst_decoder_instructionword_wire[5]), .B(imem_data[5]), 
        .S0(n504), .Y(n1228) );
  MX2X1 U1209 ( .A(inst_decoder_instructionword_wire[6]), .B(imem_data[6]), 
        .S0(n504), .Y(n1227) );
  OR2X1 U651 ( .A(pc_init[3]), .B(rstx), .Y(n965) );
  OR2X1 U624 ( .A(pc_init[4]), .B(rstx), .Y(n950) );
  OR2X1 U597 ( .A(pc_init[5]), .B(rstx), .Y(n935) );
  OR2X1 U744 ( .A(pc_init[1]), .B(rstx), .Y(n1026) );
  OR2X1 U680 ( .A(pc_init[2]), .B(rstx), .Y(n980) );
  OR2X1 U487 ( .A(pc_init[9]), .B(rstx), .Y(n875) );
  OR2X1 U570 ( .A(pc_init[6]), .B(rstx), .Y(n920) );
  OR2X1 U903 ( .A(pc_init[0]), .B(rstx), .Y(n1075) );
  OR2X1 U543 ( .A(pc_init[7]), .B(rstx), .Y(n905) );
  OR2X1 U516 ( .A(pc_init[8]), .B(rstx), .Y(n890) );
  OR2X1 U371 ( .A(pc_init[13]), .B(rstx), .Y(n815) );
  OR2X1 U458 ( .A(pc_init[10]), .B(rstx), .Y(n860) );
  OR2X1 U429 ( .A(pc_init[11]), .B(rstx), .Y(n845) );
  OR2X1 U400 ( .A(pc_init[12]), .B(rstx), .Y(n830) );
  NAND2BX1 U907 ( .AN(pc_init[14]), .B(n2261), .Y(n1078) );
  NAND2X1 U902 ( .A(pc_init[0]), .B(n2261), .Y(n1076) );
  NAND2X1 U743 ( .A(pc_init[1]), .B(n2261), .Y(n1027) );
  NAND2X1 U596 ( .A(pc_init[5]), .B(n2260), .Y(n936) );
  NAND2X1 U623 ( .A(pc_init[4]), .B(n2260), .Y(n951) );
  NAND2X1 U650 ( .A(pc_init[3]), .B(n2260), .Y(n966) );
  NAND2X1 U679 ( .A(pc_init[2]), .B(n2260), .Y(n981) );
  NAND2X1 U906 ( .A(pc_init[14]), .B(n2261), .Y(n1079) );
  AOI221X2 U156 ( .A0(ic_simm_B1_wire[24]), .A1(n2258), .B0(n2219), .B1(
        rf_RF_reg_0__24_), .C0(n136), .Y(n134) );
  AOI22X1 U88 ( .A0(n2217), .A1(rf_RF_reg_3__27_), .B0(n2215), .B1(
        rf_RF_reg_1__27_), .Y(n96) );
  AOI221X2 U86 ( .A0(ic_simm_B1_wire[27]), .A1(n2258), .B0(n2219), .B1(
        rf_RF_reg_0__27_), .C0(n94), .Y(n92) );
  AOI22X1 U25 ( .A0(n2217), .A1(rf_RF_reg_3__30_), .B0(n2215), .B1(
        rf_RF_reg_1__30_), .Y(n56) );
  AOI21X1 fu_ALU_fu_arch_U117 ( .A0(n2189), .A1(n2126), .B0(
        fu_ALU_fu_arch_n303), .Y(fu_ALU_fu_arch_n295) );
  AOI22X1 U46 ( .A0(n2217), .A1(rf_RF_reg_3__29_), .B0(n2215), .B1(
        rf_RF_reg_1__29_), .Y(n72) );
  AOI21X1 U44 ( .A0(n2220), .A1(rf_RF_reg_0__29_), .B0(n70), .Y(n68) );
  OAI21X6 fu_ALU_fu_arch_U475 ( .A0(n1769), .A1(n1774), .B0(
        fu_ALU_fu_arch_n675), .Y(fu_ALU_fu_arch_n434) );
  AOI22X1 U110 ( .A0(n2217), .A1(rf_RF_reg_3__26_), .B0(n2215), .B1(
        rf_RF_reg_1__26_), .Y(n109) );
  AOI221X2 U108 ( .A0(ic_simm_B1_wire[26]), .A1(n2258), .B0(n2219), .B1(
        rf_RF_reg_0__26_), .C0(n107), .Y(n105) );
  AOI221X2 U198 ( .A0(ic_simm_B1_wire[22]), .A1(n2258), .B0(n2219), .B1(
        rf_RF_reg_0__22_), .C0(n161), .Y(n159) );
  AOI221X2 U130 ( .A0(ic_simm_B1_wire[25]), .A1(n2258), .B0(n2219), .B1(
        rf_RF_reg_0__25_), .C0(n120), .Y(n118) );
  AOI221X2 U219 ( .A0(ic_simm_B1_wire[21]), .A1(n2258), .B0(n2219), .B1(
        rf_RF_reg_0__21_), .C0(n173), .Y(n171) );
  AOI221X2 U261 ( .A0(ic_simm_B1_wire[19]), .A1(n2258), .B0(n2219), .B1(
        rf_RF_reg_0__19_), .C0(n197), .Y(n195) );
  AOI221X2 U283 ( .A0(ic_simm_B1_wire[18]), .A1(n2258), .B0(n2219), .B1(
        rf_RF_reg_0__18_), .C0(n211), .Y(n209) );
  AOI221X2 U305 ( .A0(ic_simm_B1_wire[17]), .A1(n2258), .B0(n2219), .B1(
        rf_RF_reg_0__17_), .C0(n224), .Y(n222) );
  AOI32X2 fu_ALU_fu_arch_U385 ( .A0(n2152), .A1(fu_ALU_fu_arch_n617), .A2(
        n1762), .B0(fu_ALU_fu_arch_N628), .B1(n2192), .Y(fu_ALU_fu_arch_n615)
         );
  AOI22X2 fu_ALU_fu_arch_U384 ( .A0(n2190), .A1(n2152), .B0(n2193), .B1(
        fu_ALU_fu_arch_N49), .Y(fu_ALU_fu_arch_n616) );
  AOI221X2 U352 ( .A0(ic_simm_B1_wire[15]), .A1(n2258), .B0(n2219), .B1(
        rf_RF_reg_0__15_), .C0(n257), .Y(n255) );
  AOI22X2 fu_ALU_fu_arch_U400 ( .A0(n2154), .A1(n2190), .B0(n2193), .B1(
        fu_ALU_fu_arch_N48), .Y(fu_ALU_fu_arch_n630) );
  AOI22X1 U927 ( .A0(n2220), .A1(rf_RF_reg_0__14_), .B0(n2215), .B1(
        rf_RF_reg_1__14_), .Y(n508) );
  OAI31X4 fu_ALU_fu_arch_U485 ( .A0(fu_ALU_o1reg[12]), .A1(n2196), .A2(n1744), 
        .B0(fu_ALU_fu_arch_n685), .Y(fu_ALU_fu_arch_n679) );
  AOI22X1 U448 ( .A0(n2220), .A1(rf_RF_reg_0__11_), .B0(n2216), .B1(
        rf_RF_reg_1__11_), .Y(n301) );
  OAI211X2 fu_ALU_fu_arch_U15 ( .A0(fu_ALU_fu_arch_n125), .A1(n1745), .B0(
        fu_ALU_fu_arch_n126), .C0(fu_ALU_fu_arch_n127), .Y(fu_ALU_fu_arch_n115) );
  OAI211X2 fu_ALU_fu_arch_U34 ( .A0(fu_ALU_fu_arch_n125), .A1(n1742), .B0(
        fu_ALU_fu_arch_n151), .C0(fu_ALU_fu_arch_n152), .Y(fu_ALU_fu_arch_n145) );
  AOI22X1 U589 ( .A0(n2220), .A1(rf_RF_reg_0__6_), .B0(n2216), .B1(
        rf_RF_reg_1__6_), .Y(n359) );
  AOI22X1 U643 ( .A0(n2220), .A1(rf_RF_reg_0__4_), .B0(n2216), .B1(
        rf_RF_reg_1__4_), .Y(n379) );
  AOI22X1 U670 ( .A0(n2220), .A1(rf_RF_reg_0__3_), .B0(n2215), .B1(
        rf_RF_reg_1__3_), .Y(n389) );
  OAI31X4 fu_ALU_fu_arch_U613 ( .A0(fu_ALU_o1reg[0]), .A1(n1749), .A2(n2195), 
        .B0(fu_ALU_fu_arch_n750), .Y(fu_ALU_fu_arch_n748) );
  AOI211X4 fu_ALU_fu_arch_U612 ( .A0(n2191), .A1(fu_ALU_fu_arch_N612), .B0(
        fu_ALU_fu_arch_n747), .C0(fu_ALU_fu_arch_n748), .Y(fu_ALU_fu_arch_n742) );
  AOI21X1 U941 ( .A0(n2220), .A1(rf_RF_reg_0__31_), .B0(n516), .Y(n515) );
  NOR2X4 U1143 ( .A(n561), .B(rf_BOOL_t1opcode_wire_0_), .Y(n601) );
  AOI31X1 U1139 ( .A0(n602), .A1(n603), .A2(n559), .B0(
        inst_decoder_instructionword_wire[41]), .Y(n595) );
  OAI2BB1X1 U1018 ( .A0N(rf_RF_t1load_wire), .A1N(n2211), .B0(n550), .Y(n1131)
         );
  OAI22X1 U1026 ( .A0(n2210), .A1(n132), .B0(n544), .B1(n552), .Y(n1133) );
  AOI32X1 U1128 ( .A0(n590), .A1(n578), .A2(
        inst_decoder_instructionword_wire[36]), .B0(n2256), .B1(n2211), .Y(
        n592) );
  OAI21X1 U114 ( .A0(n112), .A1(n25), .B0(n113), .Y(n701) );
  OAI21X1 U112 ( .A0(n2254), .A1(n110), .B0(n111), .Y(n700) );
  AOI22X1 U1022 ( .A0(n2245), .A1(n220), .B0(n231), .B1(n419), .Y(n1132) );
  AOI2BB2X1 U1000 ( .B0(n2241), .B1(n220), .A0N(rf_RF_reg_0__0_), .A1N(n2242), 
        .Y(n1123) );
  OAI21X1 U134 ( .A0(n2254), .A1(n123), .B0(n124), .Y(n710) );
  OAI21X1 U160 ( .A0(n2254), .A1(n139), .B0(n140), .Y(n720) );
  OAI21X1 U181 ( .A0(n2254), .A1(n153), .B0(n154), .Y(n730) );
  AOI2BB2X1 U1006 ( .B0(n2229), .B1(n220), .A0N(rf_RF_reg_3__0_), .A1N(n2230), 
        .Y(n1126) );
  AOI2BB2X1 U1004 ( .B0(n2233), .B1(n220), .A0N(rf_RF_reg_2__0_), .A1N(n2234), 
        .Y(n1125) );
  AOI2BB2X1 U1002 ( .B0(n2237), .B1(n220), .A0N(rf_RF_reg_1__0_), .A1N(n2238), 
        .Y(n1124) );
  OAI21X1 U202 ( .A0(n2254), .A1(n165), .B0(n166), .Y(n740) );
  AOI21X1 U882 ( .A0(fu_LSU_status_addr_reg_1__3_), .A1(
        fu_LSU_status_addr_reg_1__4_), .B0(n2211), .Y(n497) );
  OAI21X1 U223 ( .A0(n2254), .A1(n177), .B0(n178), .Y(n750) );
  AOI22X1 U948 ( .A0(fu_ALU_o1reg[0]), .A1(n2252), .B0(n2251), .B1(n2111), .Y(
        n520) );
  OAI21X1 U244 ( .A0(n2254), .A1(n189), .B0(n190), .Y(n760) );
  OAI21X1 U265 ( .A0(n2255), .A1(n201), .B0(n202), .Y(n770) );
  OAI21X1 U287 ( .A0(n2255), .A1(n215), .B0(n216), .Y(n780) );
  OAI21X1 U384 ( .A0(n272), .A1(n264), .B0(n277), .Y(n827) );
  AOI22X1 U357 ( .A0(fu_ALU_fu_arch_sub_200_B_14_), .A1(n2253), .B0(n2251), 
        .B1(rf_RF_t1data_wire[14]), .Y(n261) );
  OAI21X1 U356 ( .A0(n2255), .A1(n260), .B0(n261), .Y(n810) );
  OAI21X1 U413 ( .A0(n286), .A1(n264), .B0(n288), .Y(n842) );
  AOI22X1 U365 ( .A0(fu_ALU_o1reg[13]), .A1(n2253), .B0(n2251), .B1(n1823), 
        .Y(n269) );
  OAI21X1 U364 ( .A0(n2255), .A1(n268), .B0(n269), .Y(n813) );
  OAI21X1 U309 ( .A0(n2255), .A1(n228), .B0(n229), .Y(n790) );
  AOI22X1 U394 ( .A0(fu_ALU_o1reg[12]), .A1(n2253), .B0(n2251), .B1(n1820), 
        .Y(n284) );
  OAI21X1 U393 ( .A0(n2255), .A1(n283), .B0(n284), .Y(n828) );
  AOI22X1 U335 ( .A0(n2153), .A1(n2253), .B0(n2251), .B1(rf_RF_t1data_wire[15]), .Y(n249) );
  OAI21X1 U334 ( .A0(n2255), .A1(n248), .B0(n249), .Y(n800) );
  OAI21X1 U422 ( .A0(n2255), .A1(n294), .B0(n295), .Y(n843) );
  AOI22X1 U510 ( .A0(fu_ALU_fu_arch_sub_200_B_8_), .A1(n2252), .B0(n2251), 
        .B1(rf_RF_t1data_wire[8]), .Y(n330) );
  MX2X1 U1246 ( .A(inst_fetch_N76), .B(inst_fetch_reset_cntr_30_), .S0(n2205), 
        .Y(n1264) );
  MX2X1 U1245 ( .A(inst_fetch_N75), .B(inst_fetch_reset_cntr_29_), .S0(n2204), 
        .Y(n1263) );
  MX2X1 U1216 ( .A(inst_fetch_N74), .B(inst_fetch_reset_cntr_28_), .S0(n2204), 
        .Y(n1234) );
  MX2X1 U1244 ( .A(inst_fetch_N73), .B(inst_fetch_reset_cntr_27_), .S0(n2205), 
        .Y(n1262) );
  MX2X1 U1217 ( .A(inst_fetch_N72), .B(inst_fetch_reset_cntr_26_), .S0(n2204), 
        .Y(n1235) );
  MX2X1 U1243 ( .A(inst_fetch_N71), .B(inst_fetch_reset_cntr_25_), .S0(n2204), 
        .Y(n1261) );
  OAI21X1 fu_ALU_fu_arch_U664 ( .A0(n1776), .A1(n2134), .B0(
        fu_ALU_fu_arch_n370), .Y(fu_ALU_fu_arch_n764) );
  AOI21X1 fu_ALU_fu_arch_U168 ( .A0(fu_ALU_fu_arch_n242), .A1(
        fu_ALU_fu_arch_n384), .B0(fu_ALU_fu_arch_n296), .Y(fu_ALU_fu_arch_n383) );
  AOI21X1 U23 ( .A0(n2220), .A1(rf_RF_reg_0__30_), .B0(n54), .Y(n50) );
  OAI22X1 fu_ALU_fu_arch_U120 ( .A0(n2172), .A1(fu_ALU_fu_arch_n306), .B0(
        fu_ALU_fu_arch_n307), .B1(fu_ALU_fu_arch_n308), .Y(fu_ALU_fu_arch_n305) );
  OAI22X1 fu_ALU_fu_arch_U118 ( .A0(fu_ALU_opc1reg[3]), .A1(n2188), .B0(n2126), 
        .B1(fu_ALU_opc1reg[2]), .Y(fu_ALU_fu_arch_n303) );
  AOI21X1 fu_ALU_fu_arch_U181 ( .A0(fu_ALU_fu_arch_n242), .A1(
        fu_ALU_fu_arch_n405), .B0(fu_ALU_fu_arch_n296), .Y(fu_ALU_fu_arch_n404) );
  AO21X2 fu_ALU_fu_arch_U350 ( .A0(fu_ALU_fu_arch_n590), .A1(n2105), .B0(
        fu_ALU_fu_arch_n591), .Y(fu_ALU_fu_arch_n328) );
  AOI21X4 fu_ALU_fu_arch_U372 ( .A0(n2105), .A1(fu_ALU_fu_arch_n438), .B0(
        fu_ALU_fu_arch_n606), .Y(fu_ALU_fu_arch_n536) );
  AO21X2 fu_ALU_fu_arch_U368 ( .A0(fu_ALU_fu_arch_n434), .A1(n2105), .B0(
        fu_ALU_fu_arch_n606), .Y(fu_ALU_fu_arch_n539) );
  OAI22X1 fu_ALU_fu_arch_U453 ( .A0(fu_ALU_fu_arch_n135), .A1(
        fu_ALU_fu_arch_n132), .B0(fu_ALU_fu_arch_n131), .B1(
        fu_ALU_fu_arch_n134), .Y(fu_ALU_fu_arch_n660) );
  AOI22X1 U418 ( .A0(n2214), .A1(rf_RF_reg_2__12_), .B0(n2217), .B1(
        rf_RF_reg_3__12_), .Y(n291) );
  AOI22X1 U447 ( .A0(n2214), .A1(rf_RF_reg_2__11_), .B0(n2217), .B1(
        rf_RF_reg_3__11_), .Y(n302) );
  AOI22X1 U476 ( .A0(n1777), .A1(rf_RF_reg_2__10_), .B0(n2217), .B1(
        rf_RF_reg_3__10_), .Y(n313) );
  AOI22X2 fu_ALU_fu_arch_U17 ( .A0(n2191), .A1(fu_ALU_fu_arch_N621), .B0(n2193), .B1(fu_ALU_fu_arch_N42), .Y(fu_ALU_fu_arch_n126) );
  AOI22X1 U505 ( .A0(n1777), .A1(rf_RF_reg_2__9_), .B0(n2217), .B1(
        rf_RF_reg_3__9_), .Y(n326) );
  AOI22X1 U534 ( .A0(n1777), .A1(rf_RF_reg_2__8_), .B0(n2217), .B1(
        rf_RF_reg_3__8_), .Y(n339) );
  AOI22X1 U561 ( .A0(n1777), .A1(rf_RF_reg_2__7_), .B0(n2217), .B1(
        rf_RF_reg_3__7_), .Y(n350) );
  NAND4X2 fu_ALU_fu_arch_U52 ( .A(fu_ALU_fu_arch_n180), .B(fu_ALU_fu_arch_n181), .C(fu_ALU_fu_arch_n182), .D(fu_ALU_fu_arch_n183), .Y(
        ic_socket_ALU_o1_data0_wire[6]) );
  AOI22X1 U588 ( .A0(n1777), .A1(rf_RF_reg_2__6_), .B0(n2217), .B1(
        rf_RF_reg_3__6_), .Y(n360) );
  OAI21X1 fu_ALU_fu_arch_U125 ( .A0(fu_ALU_fu_arch_n242), .A1(
        fu_ALU_fu_arch_n240), .B0(fu_ALU_fu_arch_n319), .Y(fu_ALU_fu_arch_n318) );
  NOR2X1 fu_ALU_fu_arch_U615 ( .A(fu_ALU_opc1reg[3]), .B(fu_ALU_opc1reg[1]), 
        .Y(fu_ALU_fu_arch_n751) );
  AOI221X2 U1154 ( .A0(n2258), .A1(ic_simm_B1_wire[0]), .B0(n2221), .B1(
        rf_RF_reg_4__0_), .C0(n611), .Y(n608) );
  AOI22X1 U1153 ( .A0(n2217), .A1(rf_RF_reg_3__0_), .B0(n2215), .B1(
        rf_RF_reg_1__0_), .Y(n609) );
  AOI2BB2X1 U1082 ( .B0(n2207), .B1(n575), .A0N(ic_simm_B1_wire[2]), .A1N(
        n2207), .Y(n1161) );
  AOI2BB2X1 U1083 ( .B0(n2207), .B1(n576), .A0N(ic_simm_B1_wire[0]), .A1N(
        n2207), .Y(n1162) );
  OAI21X1 U27 ( .A0(n2254), .A1(n60), .B0(n61), .Y(n660) );
  OAI21X1 U6 ( .A0(n2254), .A1(n33), .B0(n34), .Y(n650) );
  OAI21X1 U1 ( .A0(n2254), .A1(n20), .B0(n21), .Y(n648) );
  OAI21X1 U48 ( .A0(n2254), .A1(n73), .B0(n74), .Y(n670) );
  AOI32X1 U291 ( .A0(fu_LSU_o1shadow_reg_1_), .A1(n1788), .A2(n2121), .B0(
        n2123), .B1(rf_RF_t1data_wire[17]), .Y(n217) );
  AOI22X1 U70 ( .A0(fu_ALU_fu_arch_sub_200_B_27_), .A1(n2252), .B0(n2250), 
        .B1(rf_RF_t1data_wire[27]), .Y(n86) );
  OAI21X1 U69 ( .A0(n2254), .A1(n85), .B0(n86), .Y(n680) );
  AOI22X1 U91 ( .A0(n2132), .A1(n2252), .B0(n2250), .B1(rf_RF_t1data_wire[26]), 
        .Y(n98) );
  OAI21X1 U90 ( .A0(n2254), .A1(n97), .B0(n98), .Y(n690) );
  AOI22X1 U113 ( .A0(n1780), .A1(n2252), .B0(n2250), .B1(rf_RF_t1data_wire[25]), .Y(n111) );
  AOI22X1 U135 ( .A0(n2136), .A1(n2252), .B0(n2250), .B1(rf_RF_t1data_wire[24]), .Y(n124) );
  AOI22X1 U161 ( .A0(n2138), .A1(n2252), .B0(n2250), .B1(rf_RF_t1data_wire[23]), .Y(n140) );
  AOI22X1 U182 ( .A0(fu_ALU_fu_arch_sub_200_B_22_), .A1(n2252), .B0(n2250), 
        .B1(rf_RF_t1data_wire[22]), .Y(n154) );
  AOI22X1 U203 ( .A0(fu_ALU_fu_arch_sub_200_B_21_), .A1(n2252), .B0(n2250), 
        .B1(rf_RF_t1data_wire[21]), .Y(n166) );
  AOI22X1 U224 ( .A0(n2144), .A1(n2253), .B0(n2250), .B1(rf_RF_t1data_wire[20]), .Y(n178) );
  AOI22X1 U245 ( .A0(fu_ALU_fu_arch_sub_200_B_19_), .A1(n2253), .B0(n2250), 
        .B1(rf_RF_t1data_wire[19]), .Y(n190) );
  AOI22X1 U266 ( .A0(fu_ALU_fu_arch_sub_200_B_18_), .A1(n2253), .B0(n2251), 
        .B1(rf_RF_t1data_wire[18]), .Y(n202) );
  AOI22X1 U288 ( .A0(fu_ALU_o1reg[17]), .A1(n2252), .B0(n2251), .B1(
        rf_RF_t1data_wire[17]), .Y(n216) );
  AOI22X1 U310 ( .A0(fu_ALU_o1reg[16]), .A1(n2253), .B0(n2251), .B1(
        rf_RF_t1data_wire[16]), .Y(n229) );
  NOR2X4 fu_ALU_fu_arch_U662 ( .A(n2176), .B(n1768), .Y(fu_ALU_fu_arch_n248)
         );
  NAND2X5 fu_ALU_fu_arch_U370 ( .A(fu_ALU_fu_arch_n220), .B(n1851), .Y(
        fu_ALU_fu_arch_n430) );
  OAI22X1 fu_ALU_fu_arch_U677 ( .A0(fu_ALU_fu_arch_n156), .A1(n2203), .B0(
        fu_ALU_fu_arch_n154), .B1(n2106), .Y(fu_ALU_fu_arch_n762) );
  NAND2X6 fu_ALU_fu_arch_U569 ( .A(n2172), .B(n1851), .Y(fu_ALU_fu_arch_n118)
         );
  INVX5 fu_ALU_fu_arch_U568 ( .A(fu_ALU_fu_arch_n118), .Y(fu_ALU_fu_arch_n178)
         );
  NAND3X2 fu_ALU_fu_arch_U42 ( .A(fu_ALU_fu_arch_n158), .B(fu_ALU_fu_arch_n159), .C(fu_ALU_fu_arch_n160), .Y(ic_socket_ALU_o1_data0_wire[7]) );
  OAI22X1 fu_ALU_fu_arch_U621 ( .A0(fu_ALU_fu_arch_n155), .A1(
        fu_ALU_fu_arch_n544), .B0(fu_ALU_fu_arch_n157), .B1(
        fu_ALU_fu_arch_n468), .Y(fu_ALU_fu_arch_n754) );
  NAND4X4 U1151 ( .A(n607), .B(n608), .C(n609), .D(n610), .Y(
        rf_RF_t1data_wire[0]) );
  NAND2X6 fu_ALU_fu_arch_U609 ( .A(fu_ALU_fu_arch_n631), .B(n2092), .Y(
        fu_ALU_fu_arch_n153) );
  OAI211X2 fu_ALU_fu_arch_U644 ( .A0(n2189), .A1(n1749), .B0(
        fu_ALU_fu_arch_n759), .C0(n2092), .Y(fu_ALU_fu_arch_n739) );
  INVX6 fu_ALU_fu_arch_U669 ( .A(n2105), .Y(fu_ALU_fu_arch_n544) );
  AOI221X4 U671 ( .A0(n2186), .A1(ic_socket_gcu_o1_data0_wire[3]), .B0(n2257), 
        .B1(ic_socket_ALU_o1_data0_wire[3]), .C0(n392), .Y(n388) );
  AOI22X1 fu_ALU_fu_arch_U605 ( .A0(n1779), .A1(fu_ALU_fu_arch_n169), .B0(
        n2193), .B1(fu_ALU_fu_arch_N33), .Y(fu_ALU_fu_arch_n743) );
  AOI22X2 fu_ALU_fu_arch_U110 ( .A0(n2190), .A1(n2180), .B0(n2193), .B1(
        fu_ALU_fu_arch_N64), .Y(fu_ALU_fu_arch_n263) );
  AOI22X2 fu_ALU_fu_arch_U532 ( .A0(n2202), .A1(fu_ALU_fu_arch_sub_200_B_30_), 
        .B0(n2201), .B1(fu_ALU_fu_arch_sub_200_B_29_), .Y(fu_ALU_fu_arch_n707)
         );
  AOI22X2 fu_ALU_fu_arch_U599 ( .A0(n2201), .A1(fu_ALU_o1reg[24]), .B0(n2200), 
        .B1(n2138), .Y(fu_ALU_fu_arch_n736) );
  AOI21X3 fu_ALU_fu_arch_U131 ( .A0(n2200), .A1(n2166), .B0(
        fu_ALU_fu_arch_n325), .Y(fu_ALU_fu_arch_n195) );
  OAI32X4 fu_ALU_fu_arch_U88 ( .A0(fu_ALU_fu_arch_n240), .A1(
        fu_ALU_fu_arch_n241), .A2(fu_ALU_fu_arch_n242), .B0(
        fu_ALU_fu_arch_n243), .B1(fu_ALU_fu_arch_n241), .Y(fu_ALU_fu_arch_n230) );
  AOI211X4 fu_ALU_fu_arch_U133 ( .A0(fu_ALU_fu_arch_n178), .A1(
        fu_ALU_fu_arch_n328), .B0(fu_ALU_fu_arch_n329), .C0(
        fu_ALU_fu_arch_n330), .Y(fu_ALU_fu_arch_n317) );
  AOI221X4 U700 ( .A0(n2186), .A1(ic_socket_gcu_o1_data0_wire[2]), .B0(n2257), 
        .B1(ic_socket_ALU_o1_data0_wire[2]), .C0(n402), .Y(n398) );
  OAI211X4 fu_ALU_fu_arch_U259 ( .A0(fu_ALU_fu_arch_n499), .A1(
        fu_ALU_fu_arch_n468), .B0(fu_ALU_fu_arch_n488), .C0(
        fu_ALU_fu_arch_n500), .Y(fu_ALU_fu_arch_n190) );
  AOI22X4 fu_ALU_fu_arch_U334 ( .A0(fu_ALU_fu_arch_n482), .A1(n1775), .B0(
        fu_ALU_fu_arch_n167), .B1(fu_ALU_fu_arch_n249), .Y(fu_ALU_fu_arch_n574) );
  AOI221X4 U536 ( .A0(n2186), .A1(ic_socket_gcu_o1_data0_wire[8]), .B0(n2257), 
        .B1(ic_socket_ALU_o1_data0_wire[8]), .C0(n341), .Y(n337) );
  NOR2X6 fu_ALU_fu_arch_U608 ( .A(fu_ALU_fu_arch_n723), .B(fu_ALU_fu_arch_n153), .Y(fu_ALU_fu_arch_n208) );
  AOI32X2 fu_ALU_fu_arch_U67 ( .A0(fu_ALU_fu_arch_n208), .A1(
        fu_ALU_fu_arch_n209), .A2(fu_ALU_fu_arch_n210), .B0(n2039), .B1(
        fu_ALU_fu_arch_n209), .Y(fu_ALU_fu_arch_n202) );
  OAI211X4 fu_ALU_fu_arch_U308 ( .A0(n1754), .A1(n2199), .B0(
        fu_ALU_fu_arch_n552), .C0(fu_ALU_fu_arch_n553), .Y(fu_ALU_fu_arch_n199) );
  AOI211X4 fu_ALU_fu_arch_U79 ( .A0(n2103), .A1(n1803), .B0(
        fu_ALU_fu_arch_n225), .C0(fu_ALU_fu_arch_n226), .Y(fu_ALU_fu_arch_n215) );
  AOI22X2 fu_ALU_fu_arch_U135 ( .A0(n2176), .A1(fu_ALU_fu_arch_n169), .B0(
        fu_ALU_fu_arch_n333), .B1(fu_ALU_fu_arch_n334), .Y(fu_ALU_fu_arch_n332) );
  AOI22X2 U946 ( .A0(n2257), .A1(ic_socket_ALU_o1_data0_wire[31]), .B0(n2221), 
        .B1(rf_RF_reg_4__31_), .Y(n514) );
  OAI22X2 fu_ALU_fu_arch_U672 ( .A0(n2109), .A1(n1774), .B0(n1769), .B1(n2125), 
        .Y(fu_ALU_fu_arch_n765) );
  NOR2X2 fu_ALU_fu_arch_U670 ( .A(n1768), .B(fu_ALU_fu_arch_n335), .Y(
        fu_ALU_fu_arch_n247) );
  INVX2 fu_ALU_fu_arch_U295 ( .A(fu_ALU_fu_arch_n518), .Y(fu_ALU_fu_arch_n500)
         );
  AOI21X4 fu_ALU_fu_arch_U268 ( .A0(n2104), .A1(fu_ALU_fu_arch_n434), .B0(
        fu_ALU_fu_arch_n511), .Y(fu_ALU_fu_arch_n213) );
  OAI211X2 fu_ALU_fu_arch_U469 ( .A0(fu_ALU_fu_arch_n621), .A1(n2199), .B0(
        fu_ALU_fu_arch_n605), .C0(fu_ALU_fu_arch_n674), .Y(fu_ALU_fu_arch_n673) );
  OAI211X2 fu_ALU_fu_arch_U623 ( .A0(n1776), .A1(n1778), .B0(
        fu_ALU_fu_arch_n687), .C0(fu_ALU_fu_arch_n655), .Y(fu_ALU_fu_arch_n755) );
  AOI22X2 fu_ALU_fu_arch_U49 ( .A0(n2191), .A1(fu_ALU_fu_arch_N619), .B0(n2193), .B1(fu_ALU_fu_arch_N40), .Y(fu_ALU_fu_arch_n176) );
  OAI22X2 fu_ALU_fu_arch_U81 ( .A0(fu_ALU_fu_arch_n157), .A1(
        fu_ALU_fu_arch_n134), .B0(fu_ALU_fu_arch_n108), .B1(
        fu_ALU_fu_arch_n228), .Y(fu_ALU_fu_arch_n225) );
  OAI22X2 fu_ALU_fu_arch_U80 ( .A0(fu_ALU_fu_arch_n155), .A1(
        fu_ALU_fu_arch_n132), .B0(n1805), .B1(fu_ALU_fu_arch_n118), .Y(
        fu_ALU_fu_arch_n226) );
  OAI211X2 fu_ALU_fu_arch_U89 ( .A0(fu_ALU_fu_arch_n166), .A1(n2203), .B0(
        fu_ALU_fu_arch_n245), .C0(fu_ALU_fu_arch_n246), .Y(fu_ALU_fu_arch_n243) );
  AOI22X2 fu_ALU_fu_arch_U647 ( .A0(fu_ALU_fu_arch_n333), .A1(n2198), .B0(
        fu_ALU_fu_arch_n175), .B1(n1749), .Y(fu_ALU_fu_arch_n759) );
  AOI211X2 fu_ALU_fu_arch_U107 ( .A0(n2191), .A1(fu_ALU_fu_arch_N643), .B0(
        fu_ALU_fu_arch_n289), .C0(fu_ALU_fu_arch_n290), .Y(fu_ALU_fu_arch_n264) );
  DFFRHQX8 fu_ALU_o1reg_reg_12_ ( .D(n828), .CK(clk), .RN(rstx), .Q(
        fu_ALU_o1reg[12]) );
  ADDHX1 inst_fetch_add_113_U1_1_11 ( .A(inst_fetch_reset_cntr_11_), .B(
        inst_fetch_add_113_carry_11_), .CO(inst_fetch_add_113_carry_12_), .S(
        inst_fetch_N57) );
  ADDHX1 inst_fetch_add_113_U1_1_10 ( .A(inst_fetch_reset_cntr_10_), .B(
        inst_fetch_add_113_carry_10_), .CO(inst_fetch_add_113_carry_11_), .S(
        inst_fetch_N56) );
  ADDHX1 inst_fetch_add_113_U1_1_4 ( .A(inst_fetch_reset_cntr_4_), .B(
        inst_fetch_add_113_carry_4_), .CO(inst_fetch_add_113_carry_5_), .S(
        inst_fetch_N50) );
  ADDHX1 inst_fetch_add_113_U1_1_8 ( .A(inst_fetch_reset_cntr_8_), .B(
        inst_fetch_add_113_carry_8_), .CO(inst_fetch_add_113_carry_9_), .S(
        inst_fetch_N54) );
  ADDHX1 inst_fetch_add_113_U1_1_14 ( .A(inst_fetch_reset_cntr_14_), .B(
        inst_fetch_add_113_carry_14_), .CO(inst_fetch_add_113_carry_15_), .S(
        inst_fetch_N60) );
  ADDHX1 inst_fetch_add_113_U1_1_18 ( .A(inst_fetch_reset_cntr_18_), .B(
        inst_fetch_add_113_carry_18_), .CO(inst_fetch_add_113_carry_19_), .S(
        inst_fetch_N64) );
  ADDHX1 inst_fetch_add_113_U1_1_21 ( .A(inst_fetch_reset_cntr_21_), .B(
        inst_fetch_add_113_carry_21_), .CO(inst_fetch_add_113_carry_22_), .S(
        inst_fetch_N67) );
  ADDHX1 inst_fetch_add_113_U1_1_19 ( .A(inst_fetch_reset_cntr_19_), .B(
        inst_fetch_add_113_carry_19_), .CO(inst_fetch_add_113_carry_20_), .S(
        inst_fetch_N65) );
  ADDHX1 inst_fetch_add_113_U1_1_15 ( .A(inst_fetch_reset_cntr_15_), .B(
        inst_fetch_add_113_carry_15_), .CO(inst_fetch_add_113_carry_16_), .S(
        inst_fetch_N61) );
  ADDHX1 inst_fetch_add_113_U1_1_2 ( .A(inst_fetch_reset_cntr_2_), .B(
        inst_fetch_add_113_carry_2_), .CO(inst_fetch_add_113_carry_3_), .S(
        inst_fetch_N48) );
  ADDHX1 inst_fetch_add_113_U1_1_20 ( .A(inst_fetch_reset_cntr_20_), .B(
        inst_fetch_add_113_carry_20_), .CO(inst_fetch_add_113_carry_21_), .S(
        inst_fetch_N66) );
  ADDHX1 inst_fetch_add_113_U1_1_3 ( .A(inst_fetch_reset_cntr_3_), .B(
        inst_fetch_add_113_carry_3_), .CO(inst_fetch_add_113_carry_4_), .S(
        inst_fetch_N49) );
  ADDHX1 inst_fetch_add_113_U1_1_9 ( .A(inst_fetch_reset_cntr_9_), .B(
        inst_fetch_add_113_carry_9_), .CO(inst_fetch_add_113_carry_10_), .S(
        inst_fetch_N55) );
  ADDHX1 inst_fetch_add_113_U1_1_22 ( .A(inst_fetch_reset_cntr_22_), .B(
        inst_fetch_add_113_carry_22_), .CO(inst_fetch_add_113_carry_23_), .S(
        inst_fetch_N68) );
  ADDHX1 inst_fetch_add_113_U1_1_7 ( .A(inst_fetch_reset_cntr_7_), .B(
        inst_fetch_add_113_carry_7_), .CO(inst_fetch_add_113_carry_8_), .S(
        inst_fetch_N53) );
  ADDHX1 inst_fetch_add_113_U1_1_6 ( .A(inst_fetch_reset_cntr_6_), .B(
        inst_fetch_add_113_carry_6_), .CO(inst_fetch_add_113_carry_7_), .S(
        inst_fetch_N52) );
  ADDHX1 inst_fetch_add_113_U1_1_17 ( .A(inst_fetch_reset_cntr_17_), .B(
        inst_fetch_add_113_carry_17_), .CO(inst_fetch_add_113_carry_18_), .S(
        inst_fetch_N63) );
  ADDHX1 inst_fetch_add_113_U1_1_5 ( .A(inst_fetch_reset_cntr_5_), .B(
        inst_fetch_add_113_carry_5_), .CO(inst_fetch_add_113_carry_6_), .S(
        inst_fetch_N51) );
  ADDHX1 inst_fetch_add_113_U1_1_23 ( .A(inst_fetch_reset_cntr_23_), .B(
        inst_fetch_add_113_carry_23_), .CO(inst_fetch_add_113_carry_24_), .S(
        inst_fetch_N69) );
  ADDHX1 inst_fetch_add_113_U1_1_1 ( .A(inst_fetch_reset_cntr_1_), .B(
        inst_fetch_reset_cntr_0_), .CO(inst_fetch_add_113_carry_2_), .S(
        inst_fetch_N47) );
  ADDHX1 inst_fetch_add_113_U1_1_12 ( .A(inst_fetch_reset_cntr_12_), .B(
        inst_fetch_add_113_carry_12_), .CO(inst_fetch_add_113_carry_13_), .S(
        inst_fetch_N58) );
  ADDHX1 inst_fetch_add_113_U1_1_16 ( .A(inst_fetch_reset_cntr_16_), .B(
        inst_fetch_add_113_carry_16_), .CO(inst_fetch_add_113_carry_17_), .S(
        inst_fetch_N62) );
  ADDHX1 inst_fetch_add_113_U1_1_13 ( .A(inst_fetch_reset_cntr_13_), .B(
        inst_fetch_add_113_carry_13_), .CO(inst_fetch_add_113_carry_14_), .S(
        inst_fetch_N59) );
  ADDHX1 inst_fetch_add_113_U1_1_24 ( .A(inst_fetch_reset_cntr_24_), .B(
        inst_fetch_add_113_carry_24_), .CO(inst_fetch_add_113_carry_25_), .S(
        inst_fetch_N70) );
  ADDHX1 inst_fetch_add_113_U1_1_25 ( .A(inst_fetch_reset_cntr_25_), .B(
        inst_fetch_add_113_carry_25_), .CO(inst_fetch_add_113_carry_26_), .S(
        inst_fetch_N71) );
  ADDHX1 inst_fetch_add_113_U1_1_26 ( .A(inst_fetch_reset_cntr_26_), .B(
        inst_fetch_add_113_carry_26_), .CO(inst_fetch_add_113_carry_27_), .S(
        inst_fetch_N72) );
  ADDHX1 inst_fetch_add_113_U1_1_27 ( .A(inst_fetch_reset_cntr_27_), .B(
        inst_fetch_add_113_carry_27_), .CO(inst_fetch_add_113_carry_28_), .S(
        inst_fetch_N73) );
  ADDHX1 inst_fetch_add_113_U1_1_30 ( .A(inst_fetch_reset_cntr_30_), .B(
        inst_fetch_add_113_carry_30_), .CO(inst_fetch_add_113_carry_31_), .S(
        inst_fetch_N76) );
  ADDHX1 inst_fetch_add_113_U1_1_29 ( .A(inst_fetch_reset_cntr_29_), .B(
        inst_fetch_add_113_carry_29_), .CO(inst_fetch_add_113_carry_30_), .S(
        inst_fetch_N75) );
  ADDHX1 inst_fetch_add_113_U1_1_28 ( .A(inst_fetch_reset_cntr_28_), .B(
        inst_fetch_add_113_carry_28_), .CO(inst_fetch_add_113_carry_29_), .S(
        inst_fetch_N74) );
  ADDFX1 fu_ALU_fu_arch_sub_200_U2_31 ( .A(n2180), .B(n1774), .CI(
        fu_ALU_fu_arch_sub_200_carry_31_), .S(fu_ALU_fu_arch_N643) );
  ADDFX1 fu_ALU_fu_arch_sub_200_U2_1 ( .A(fu_ALU_fu_arch_sub_200_A_1_), .B(
        n1738), .CI(fu_ALU_fu_arch_sub_200_carry_1_), .CO(
        fu_ALU_fu_arch_sub_200_carry_2_), .S(fu_ALU_fu_arch_N613) );
  ADDFX1 fu_ALU_fu_arch_sub_200_U2_2 ( .A(n2176), .B(
        fu_ALU_fu_arch_sub_200_B_not_2_), .CI(fu_ALU_fu_arch_sub_200_carry_2_), 
        .CO(fu_ALU_fu_arch_sub_200_carry_3_), .S(fu_ALU_fu_arch_N614) );
  ADDFX1 fu_ALU_fu_arch_sub_200_U2_3 ( .A(n2174), .B(n1773), .CI(
        fu_ALU_fu_arch_sub_200_carry_3_), .CO(fu_ALU_fu_arch_sub_200_carry_4_), 
        .S(fu_ALU_fu_arch_N615) );
  ADDFX1 fu_ALU_fu_arch_sub_200_U2_4 ( .A(n2172), .B(
        fu_ALU_fu_arch_sub_200_B_not_4_), .CI(fu_ALU_fu_arch_sub_200_carry_4_), 
        .CO(fu_ALU_fu_arch_sub_200_carry_5_), .S(fu_ALU_fu_arch_N616) );
  ADDFX1 fu_ALU_fu_arch_sub_200_U2_5 ( .A(fu_ALU_t1reg[5]), .B(n1754), .CI(
        fu_ALU_fu_arch_sub_200_carry_5_), .CO(fu_ALU_fu_arch_sub_200_carry_6_), 
        .S(fu_ALU_fu_arch_N617) );
  ADDFX1 fu_ALU_fu_arch_sub_200_U2_6 ( .A(n2169), .B(
        fu_ALU_fu_arch_sub_200_B_not_6_), .CI(fu_ALU_fu_arch_sub_200_carry_6_), 
        .CO(fu_ALU_fu_arch_sub_200_carry_7_), .S(fu_ALU_fu_arch_N618) );
  ADDFX1 fu_ALU_fu_arch_sub_200_U2_7 ( .A(n2167), .B(n1743), .CI(
        fu_ALU_fu_arch_sub_200_carry_7_), .CO(fu_ALU_fu_arch_sub_200_carry_8_), 
        .S(fu_ALU_fu_arch_N619) );
  ADDFX1 fu_ALU_fu_arch_sub_200_U2_8 ( .A(n2165), .B(n2164), .CI(
        fu_ALU_fu_arch_sub_200_carry_8_), .CO(fu_ALU_fu_arch_sub_200_carry_9_), 
        .S(fu_ALU_fu_arch_N620) );
  ADDFX1 fu_ALU_fu_arch_add_171_U1_1 ( .A(fu_ALU_fu_arch_sub_200_A_1_), .B(
        n2177), .CI(fu_ALU_fu_arch_add_171_carry_1_), .CO(
        fu_ALU_fu_arch_add_171_carry_2_), .S(fu_ALU_fu_arch_N34) );
  ADDFX1 fu_ALU_fu_arch_add_171_U1_2 ( .A(n2176), .B(
        fu_ALU_fu_arch_sub_200_B_2_), .CI(fu_ALU_fu_arch_add_171_carry_2_), 
        .CO(fu_ALU_fu_arch_add_171_carry_3_), .S(fu_ALU_fu_arch_N35) );
  ADDFX1 fu_ALU_fu_arch_add_171_U1_3 ( .A(n2174), .B(n2173), .CI(
        fu_ALU_fu_arch_add_171_carry_3_), .CO(fu_ALU_fu_arch_add_171_carry_4_), 
        .S(fu_ALU_fu_arch_N36) );
  ADDFX1 fu_ALU_fu_arch_add_171_U1_4 ( .A(n2172), .B(
        fu_ALU_fu_arch_sub_200_B_4_), .CI(fu_ALU_fu_arch_add_171_carry_4_), 
        .CO(fu_ALU_fu_arch_add_171_carry_5_), .S(fu_ALU_fu_arch_N37) );
  ADDFX1 fu_ALU_fu_arch_add_171_U1_5 ( .A(fu_ALU_t1reg[5]), .B(
        fu_ALU_fu_arch_sub_200_B_5_), .CI(fu_ALU_fu_arch_add_171_carry_5_), 
        .CO(fu_ALU_fu_arch_add_171_carry_6_), .S(fu_ALU_fu_arch_N38) );
  ADDFX1 fu_ALU_fu_arch_add_171_U1_6 ( .A(n2169), .B(n2168), .CI(
        fu_ALU_fu_arch_add_171_carry_6_), .CO(fu_ALU_fu_arch_add_171_carry_7_), 
        .S(fu_ALU_fu_arch_N39) );
  ADDFX1 fu_ALU_fu_arch_add_171_U1_7 ( .A(n2167), .B(n2166), .CI(
        fu_ALU_fu_arch_add_171_carry_7_), .CO(fu_ALU_fu_arch_add_171_carry_8_), 
        .S(fu_ALU_fu_arch_N40) );
  ADDFX1 fu_ALU_fu_arch_add_171_U1_8 ( .A(n2165), .B(
        fu_ALU_fu_arch_sub_200_B_8_), .CI(fu_ALU_fu_arch_add_171_carry_8_), 
        .CO(fu_ALU_fu_arch_add_171_carry_9_), .S(fu_ALU_fu_arch_N41) );
  ADDFX1 fu_ALU_fu_arch_add_171_U1_9 ( .A(n2163), .B(
        fu_ALU_fu_arch_sub_200_B_9_), .CI(fu_ALU_fu_arch_add_171_carry_9_), 
        .CO(fu_ALU_fu_arch_add_171_carry_10_), .S(fu_ALU_fu_arch_N42) );
  ADDFX1 fu_ALU_fu_arch_add_171_U1_31 ( .A(n2180), .B(n2124), .CI(
        fu_ALU_fu_arch_add_171_carry_31_), .S(fu_ALU_fu_arch_N64) );
  DFFRHQX8 fu_ALU_opc1reg_reg_3_ ( .D(n1119), .CK(clk), .RN(rstx), .Q(
        fu_ALU_opc1reg[3]) );
  DFFRHQX8 fu_ALU_o1reg_reg_17_ ( .D(n780), .CK(clk), .RN(rstx), .Q(
        fu_ALU_o1reg[17]) );
  DFFRHQX8 fu_ALU_o1reg_reg_6_ ( .D(n918), .CK(clk), .RN(rstx), .Q(
        fu_ALU_o1reg[6]) );
  DFFRHQX8 inst_decoder_socket_lsu_o1_bus_cntrl_reg_reg_0_ ( .D(n1188), .CK(
        clk), .RN(rstx), .Q(ic_socket_lsu_o1_bus_cntrl_wire_0_) );
  DFFRHQX8 fu_ALU_opc1reg_reg_0_ ( .D(n1115), .CK(clk), .RN(rstx), .Q(
        fu_ALU_opc1reg[0]) );
  DFFRHQX8 fu_ALU_o1reg_reg_22_ ( .D(n730), .CK(clk), .RN(rstx), .Q(
        fu_ALU_o1reg[22]) );
  DFFRHQX8 fu_ALU_o1reg_reg_20_ ( .D(n750), .CK(clk), .RN(rstx), .Q(
        fu_ALU_o1reg[20]) );
  DFFRHQX8 fu_ALU_o1reg_reg_31_ ( .D(n648), .CK(clk), .RN(rstx), .Q(
        fu_ALU_o1reg[31]) );
  DFFRHQX8 fu_ALU_o1reg_reg_23_ ( .D(n720), .CK(clk), .RN(rstx), .Q(
        fu_ALU_o1reg[23]) );
  DFFRHQX8 fu_LSU_status_addr_reg_reg_1__3_ ( .D(n1107), .CK(clk), .RN(rstx), 
        .Q(fu_LSU_status_addr_reg_1__3_) );
  DFFRHQX8 fu_ALU_o1reg_reg_13_ ( .D(n813), .CK(clk), .RN(rstx), .Q(
        fu_ALU_o1reg[13]) );
  DFFRQX4 inst_fetch_instruction_reg_reg_37_ ( .D(n1196), .CK(clk), .RN(rstx), 
        .Q(inst_decoder_instructionword_wire[37]) );
  DFFRQX4 inst_fetch_instruction_reg_reg_36_ ( .D(n1197), .CK(clk), .RN(rstx), 
        .Q(inst_decoder_instructionword_wire[36]) );
  DFFRHQX8 fu_ALU_o1reg_reg_10_ ( .D(n858), .CK(clk), .RN(rstx), .Q(
        fu_ALU_o1reg[10]) );
  DFFRHQX8 fu_ALU_o1reg_reg_3_ ( .D(n963), .CK(clk), .RN(rstx), .Q(
        fu_ALU_o1reg[3]) );
  DFFRQX4 fu_ALU_o1reg_reg_14_ ( .D(n810), .CK(clk), .RN(rstx), .Q(
        fu_ALU_o1reg[14]) );
  DFFRQX4 fu_ALU_o1reg_reg_29_ ( .D(n660), .CK(clk), .RN(rstx), .Q(
        fu_ALU_o1reg[29]) );
  DFFRQX4 inst_decoder_rf_RF_wr_opc_reg_reg_2_ ( .D(n1130), .CK(clk), .RN(rstx), .Q(rf_RF_t1opcode_wire[2]) );
  DFFRQX4 inst_decoder_fu_gcu_ra_load_reg_reg ( .D(n1146), .CK(clk), .RN(rstx), 
        .Q(inst_fetch_ra_load_wire) );
  DFFRQX4 inst_fetch_reset_cntr_reg_21_ ( .D(n1259), .CK(clk), .RN(rstx), .Q(
        inst_fetch_reset_cntr_21_) );
  DFFRQX4 inst_fetch_reset_cntr_reg_28_ ( .D(n1234), .CK(clk), .RN(rstx), .Q(
        inst_fetch_reset_cntr_28_) );
  DFFRQX4 inst_fetch_reset_cntr_reg_24_ ( .D(n1236), .CK(clk), .RN(rstx), .Q(
        inst_fetch_reset_cntr_24_) );
  DFFRQX4 inst_fetch_reset_cntr_reg_13_ ( .D(n1255), .CK(clk), .RN(rstx), .Q(
        inst_fetch_reset_cntr_13_) );
  DFFRQX4 inst_fetch_reset_cntr_reg_17_ ( .D(n1257), .CK(clk), .RN(rstx), .Q(
        inst_fetch_reset_cntr_17_) );
  DFFRQX4 inst_fetch_reset_cntr_reg_4_ ( .D(n1246), .CK(clk), .RN(rstx), .Q(
        inst_fetch_reset_cntr_4_) );
  DFFRQX4 inst_fetch_reset_cntr_reg_6_ ( .D(n1245), .CK(clk), .RN(rstx), .Q(
        inst_fetch_reset_cntr_6_) );
  DFFRQX4 inst_fetch_reset_cntr_reg_8_ ( .D(n1244), .CK(clk), .RN(rstx), .Q(
        inst_fetch_reset_cntr_8_) );
  DFFRQX4 inst_fetch_reset_cntr_reg_9_ ( .D(n1253), .CK(clk), .RN(rstx), .Q(
        inst_fetch_reset_cntr_9_) );
  DFFRQX4 inst_decoder_rf_RF_wr_opc_reg_reg_1_ ( .D(n1128), .CK(clk), .RN(rstx), .Q(rf_RF_t1opcode_wire[1]) );
  DFFRQX4 inst_fetch_instruction_reg_reg_39_ ( .D(n1194), .CK(clk), .RN(rstx), 
        .Q(inst_decoder_instructionword_wire[39]) );
  DFFRQX4 rf_BOOL_reg_reg_0__0_ ( .D(n1136), .CK(clk), .RN(rstx), .Q(
        rf_BOOL_reg_0__0_) );
  DFFRQX4 fu_ALU_o1reg_reg_0_ ( .D(n1098), .CK(clk), .RN(rstx), .Q(
        fu_ALU_o1reg[0]) );
  DFFSQX2 inst_fetch_reset_lock_reg ( .D(n1191), .CK(clk), .SN(rstx), .Q(
        inst_fetch_reset_lock) );
  DFFSQX2 fu_LSU_wr_en_x_reg_reg_0_ ( .D(n1099), .CK(clk), .SN(rstx), .Q(
        fu_LSU_wr_en_x[0]) );
  DFFSQX2 fu_LSU_mem_en_x_reg_reg_0_ ( .D(n1111), .CK(clk), .SN(rstx), .Q(
        fu_LSU_mem_en_x[0]) );
  DFFRQX4 inst_fetch_reset_cntr_reg_22_ ( .D(n1237), .CK(clk), .RN(rstx), .Q(
        inst_fetch_reset_cntr_22_) );
  DFFRQX4 inst_fetch_reset_cntr_reg_23_ ( .D(n1260), .CK(clk), .RN(rstx), .Q(
        inst_fetch_reset_cntr_23_) );
  DFFRHQX8 inst_fetch_instruction_reg_reg_1_ ( .D(n1232), .CK(clk), .RN(rstx), 
        .Q(inst_decoder_N121) );
  DFFRHQX8 fu_ALU_t1reg_reg_5_ ( .D(n938), .CK(clk), .RN(rstx), .Q(
        fu_ALU_t1reg[5]) );
  DFFRQX4 inst_decoder_fu_LSU_opc_reg_reg_2_ ( .D(n1110), .CK(clk), .RN(rstx), 
        .Q(fu_LSU_t1opcode_wire[2]) );
  DFFRQX4 inst_fetch_instruction_reg_reg_41_ ( .D(n1192), .CK(clk), .RN(rstx), 
        .Q(inst_decoder_instructionword_wire[41]) );
  DFFRQX4 inst_decoder_rf_BOOL_wr_opc_reg_reg_0_ ( .D(n1137), .CK(clk), .RN(
        rstx), .Q(rf_BOOL_t1opcode_wire_0_) );
  DFFRHQX8 fu_ALU_o1reg_reg_24_ ( .D(n710), .CK(clk), .RN(rstx), .Q(
        fu_ALU_o1reg[24]) );
  DFFRHQX8 fu_ALU_opc1reg_reg_1_ ( .D(n1117), .CK(clk), .RN(rstx), .Q(
        fu_ALU_opc1reg[1]) );
  DFFRHQX8 fu_ALU_opc1reg_reg_2_ ( .D(n1113), .CK(clk), .RN(rstx), .Q(
        fu_ALU_opc1reg[2]) );
  DFFRHQX8 fu_ALU_o1reg_reg_16_ ( .D(n790), .CK(clk), .RN(rstx), .Q(
        fu_ALU_o1reg[16]) );
  DFFRHQX8 inst_decoder_fu_LIFTING_opc_reg_reg_1_ ( .D(n1139), .CK(clk), .RN(
        rstx), .Q(fu_LIFTING_t1opcode_wire[1]) );
  DFFRHQX8 inst_decoder_fu_LIFTING_opc_reg_reg_2_ ( .D(n1141), .CK(clk), .RN(
        rstx), .Q(fu_LIFTING_t1opcode_wire[2]) );
  DFFRHQX8 inst_fetch_instruction_reg_reg_35_ ( .D(n1198), .CK(clk), .RN(rstx), 
        .Q(inst_decoder_instructionword_wire[35]) );
  DFFRHQX8 inst_decoder_fu_LIFTING_opc_reg_reg_0_ ( .D(n1140), .CK(clk), .RN(
        rstx), .Q(fu_LIFTING_t1opcode_wire[0]) );
  DFFRHQX8 inst_decoder_fu_LSU_opc_reg_reg_1_ ( .D(n1104), .CK(clk), .RN(rstx), 
        .Q(fu_LSU_t1opcode_wire[1]) );
  DFFRHQX8 inst_fetch_instruction_reg_reg_2_ ( .D(n1231), .CK(clk), .RN(rstx), 
        .Q(inst_decoder_N230) );
  DFFRHQX8 fu_LSU_status_addr_reg_reg_1__4_ ( .D(n1105), .CK(clk), .RN(rstx), 
        .Q(fu_LSU_status_addr_reg_1__4_) );
  DFFRHQX8 inst_fetch_instruction_reg_reg_3_ ( .D(n1230), .CK(clk), .RN(rstx), 
        .Q(inst_decoder_N232) );
  DFFRQX4 fu_ALU_o1reg_reg_25_ ( .D(n700), .CK(clk), .RN(rstx), .Q(
        fu_ALU_o1reg[25]) );
  DFFRQX4 inst_fetch_instruction_reg_reg_40_ ( .D(n1193), .CK(clk), .RN(rstx), 
        .Q(inst_decoder_instructionword_wire[40]) );
  DFFRQX4 inst_fetch_instruction_reg_reg_4_ ( .D(n1229), .CK(clk), .RN(rstx), 
        .Q(inst_decoder_instructionword_wire[4]) );
  DFFRQX4 inst_decoder_rf_RF_rd_opc_reg_reg_1_ ( .D(n1180), .CK(clk), .RN(rstx), .Q(rf_RF_r1opcode_wire[1]) );
  DFFRQX4 inst_fetch_reset_cntr_reg_20_ ( .D(n1238), .CK(clk), .RN(rstx), .Q(
        inst_fetch_reset_cntr_20_) );
  DFFRQX4 inst_fetch_reset_cntr_reg_29_ ( .D(n1263), .CK(clk), .RN(rstx), .Q(
        inst_fetch_reset_cntr_29_) );
  DFFRQX4 inst_fetch_reset_cntr_reg_25_ ( .D(n1261), .CK(clk), .RN(rstx), .Q(
        inst_fetch_reset_cntr_25_) );
  DFFRQX4 inst_fetch_reset_cntr_reg_14_ ( .D(n1241), .CK(clk), .RN(rstx), .Q(
        inst_fetch_reset_cntr_14_) );
  DFFRQX4 inst_fetch_reset_cntr_reg_18_ ( .D(n1239), .CK(clk), .RN(rstx), .Q(
        inst_fetch_reset_cntr_18_) );
  DFFRQX4 inst_fetch_reset_cntr_reg_30_ ( .D(n1264), .CK(clk), .RN(rstx), .Q(
        inst_fetch_reset_cntr_30_) );
  DFFRQX4 inst_fetch_reset_cntr_reg_27_ ( .D(n1262), .CK(clk), .RN(rstx), .Q(
        inst_fetch_reset_cntr_27_) );
  DFFRQX4 inst_fetch_reset_cntr_reg_1_ ( .D(n1249), .CK(clk), .RN(rstx), .Q(
        inst_fetch_reset_cntr_1_) );
  DFFRQX4 inst_fetch_reset_cntr_reg_16_ ( .D(n1240), .CK(clk), .RN(rstx), .Q(
        inst_fetch_reset_cntr_16_) );
  DFFRQX4 inst_fetch_reset_cntr_reg_12_ ( .D(n1242), .CK(clk), .RN(rstx), .Q(
        inst_fetch_reset_cntr_12_) );
  DFFRQX4 inst_fetch_reset_cntr_reg_7_ ( .D(n1252), .CK(clk), .RN(rstx), .Q(
        inst_fetch_reset_cntr_7_) );
  DFFRQX4 inst_fetch_reset_cntr_reg_11_ ( .D(n1254), .CK(clk), .RN(rstx), .Q(
        inst_fetch_reset_cntr_11_) );
  DFFRQX4 inst_fetch_reset_cntr_reg_2_ ( .D(n1247), .CK(clk), .RN(rstx), .Q(
        inst_fetch_reset_cntr_2_) );
  DFFRQX4 inst_fetch_reset_cntr_reg_26_ ( .D(n1235), .CK(clk), .RN(rstx), .Q(
        inst_fetch_reset_cntr_26_) );
  DFFRQX4 inst_fetch_reset_cntr_reg_15_ ( .D(n1256), .CK(clk), .RN(rstx), .Q(
        inst_fetch_reset_cntr_15_) );
  DFFRQX4 inst_fetch_reset_cntr_reg_19_ ( .D(n1258), .CK(clk), .RN(rstx), .Q(
        inst_fetch_reset_cntr_19_) );
  DFFRQX4 inst_fetch_reset_cntr_reg_3_ ( .D(n1250), .CK(clk), .RN(rstx), .Q(
        inst_fetch_reset_cntr_3_) );
  DFFRQX4 inst_fetch_reset_cntr_reg_5_ ( .D(n1251), .CK(clk), .RN(rstx), .Q(
        inst_fetch_reset_cntr_5_) );
  DFFRQX4 inst_decoder_rf_RF_wr_opc_reg_reg_0_ ( .D(n1129), .CK(clk), .RN(rstx), .Q(rf_RF_t1opcode_wire[0]) );
  DFFRQX4 inst_fetch_reset_cntr_reg_31_ ( .D(n1265), .CK(clk), .RN(rstx), .Q(
        inst_fetch_reset_cntr_31_) );
  DFFRQX4 fu_LSU_status_addr_reg_reg_1__2_ ( .D(n1100), .CK(clk), .RN(rstx), 
        .Q(fu_LSU_status_addr_reg_1__2_) );
  DFFSQX2 fu_LSU_wr_mask_x_reg_reg_0_ ( .D(n997), .CK(clk), .SN(rstx), .Q(
        fu_LSU_wr_mask_x[0]) );
  DFFSQX2 fu_LSU_wr_mask_x_reg_reg_31_ ( .D(n1025), .CK(clk), .SN(rstx), .Q(
        fu_LSU_wr_mask_x[31]) );
  DFFSQX2 fu_LSU_wr_mask_x_reg_reg_1_ ( .D(n998), .CK(clk), .SN(rstx), .Q(
        fu_LSU_wr_mask_x[1]) );
  DFFSQX2 fu_LSU_wr_mask_x_reg_reg_30_ ( .D(n1018), .CK(clk), .SN(rstx), .Q(
        fu_LSU_wr_mask_x[30]) );
  DFFSQX2 fu_LSU_wr_mask_x_reg_reg_2_ ( .D(n996), .CK(clk), .SN(rstx), .Q(
        fu_LSU_wr_mask_x[2]) );
  DFFSQX2 fu_LSU_wr_mask_x_reg_reg_29_ ( .D(n1024), .CK(clk), .SN(rstx), .Q(
        fu_LSU_wr_mask_x[29]) );
  DFFSQX2 fu_LSU_wr_mask_x_reg_reg_3_ ( .D(n999), .CK(clk), .SN(rstx), .Q(
        fu_LSU_wr_mask_x[3]) );
  DFFSQX2 fu_LSU_wr_mask_x_reg_reg_28_ ( .D(n1019), .CK(clk), .SN(rstx), .Q(
        fu_LSU_wr_mask_x[28]) );
  DFFSQX2 fu_LSU_wr_mask_x_reg_reg_4_ ( .D(n995), .CK(clk), .SN(rstx), .Q(
        fu_LSU_wr_mask_x[4]) );
  DFFSQX2 fu_LSU_wr_mask_x_reg_reg_27_ ( .D(n1023), .CK(clk), .SN(rstx), .Q(
        fu_LSU_wr_mask_x[27]) );
  DFFSQX2 fu_LSU_wr_mask_x_reg_reg_5_ ( .D(n1000), .CK(clk), .SN(rstx), .Q(
        fu_LSU_wr_mask_x[5]) );
  DFFSQX2 fu_LSU_wr_mask_x_reg_reg_26_ ( .D(n1020), .CK(clk), .SN(rstx), .Q(
        fu_LSU_wr_mask_x[26]) );
  DFFSQX2 fu_LSU_wr_mask_x_reg_reg_6_ ( .D(n994), .CK(clk), .SN(rstx), .Q(
        fu_LSU_wr_mask_x[6]) );
  DFFSQX2 fu_LSU_wr_mask_x_reg_reg_25_ ( .D(n1022), .CK(clk), .SN(rstx), .Q(
        fu_LSU_wr_mask_x[25]) );
  DFFSQX2 fu_LSU_wr_mask_x_reg_reg_7_ ( .D(n1001), .CK(clk), .SN(rstx), .Q(
        fu_LSU_wr_mask_x[7]) );
  DFFSQX2 fu_LSU_wr_mask_x_reg_reg_24_ ( .D(n1021), .CK(clk), .SN(rstx), .Q(
        fu_LSU_wr_mask_x[24]) );
  DFFSQX2 fu_LSU_wr_mask_x_reg_reg_8_ ( .D(n1005), .CK(clk), .SN(rstx), .Q(
        fu_LSU_wr_mask_x[8]) );
  DFFSQX2 fu_LSU_wr_mask_x_reg_reg_23_ ( .D(n1017), .CK(clk), .SN(rstx), .Q(
        fu_LSU_wr_mask_x[23]) );
  DFFSQX2 fu_LSU_wr_mask_x_reg_reg_9_ ( .D(n1006), .CK(clk), .SN(rstx), .Q(
        fu_LSU_wr_mask_x[9]) );
  DFFSQX2 fu_LSU_wr_mask_x_reg_reg_22_ ( .D(n1010), .CK(clk), .SN(rstx), .Q(
        fu_LSU_wr_mask_x[22]) );
  DFFSQX2 fu_LSU_wr_mask_x_reg_reg_10_ ( .D(n1004), .CK(clk), .SN(rstx), .Q(
        fu_LSU_wr_mask_x[10]) );
  DFFSQX2 fu_LSU_wr_mask_x_reg_reg_21_ ( .D(n1016), .CK(clk), .SN(rstx), .Q(
        fu_LSU_wr_mask_x[21]) );
  DFFSQX2 fu_LSU_wr_mask_x_reg_reg_11_ ( .D(n1007), .CK(clk), .SN(rstx), .Q(
        fu_LSU_wr_mask_x[11]) );
  DFFSQX2 fu_LSU_wr_mask_x_reg_reg_20_ ( .D(n1011), .CK(clk), .SN(rstx), .Q(
        fu_LSU_wr_mask_x[20]) );
  DFFSQX2 fu_LSU_wr_mask_x_reg_reg_12_ ( .D(n1003), .CK(clk), .SN(rstx), .Q(
        fu_LSU_wr_mask_x[12]) );
  DFFSQX2 fu_LSU_wr_mask_x_reg_reg_19_ ( .D(n1015), .CK(clk), .SN(rstx), .Q(
        fu_LSU_wr_mask_x[19]) );
  DFFSQX2 fu_LSU_wr_mask_x_reg_reg_13_ ( .D(n1008), .CK(clk), .SN(rstx), .Q(
        fu_LSU_wr_mask_x[13]) );
  DFFSQX2 fu_LSU_wr_mask_x_reg_reg_18_ ( .D(n1012), .CK(clk), .SN(rstx), .Q(
        fu_LSU_wr_mask_x[18]) );
  DFFSQX2 fu_LSU_wr_mask_x_reg_reg_14_ ( .D(n1002), .CK(clk), .SN(rstx), .Q(
        fu_LSU_wr_mask_x[14]) );
  DFFSQX2 fu_LSU_wr_mask_x_reg_reg_17_ ( .D(n1014), .CK(clk), .SN(rstx), .Q(
        fu_LSU_wr_mask_x[17]) );
  DFFSQX2 fu_LSU_wr_mask_x_reg_reg_15_ ( .D(n1009), .CK(clk), .SN(rstx), .Q(
        fu_LSU_wr_mask_x[15]) );
  DFFSQX2 fu_LSU_wr_mask_x_reg_reg_16_ ( .D(n1013), .CK(clk), .SN(rstx), .Q(
        fu_LSU_wr_mask_x[16]) );
  DFFRQX4 fu_ALU_o1reg_reg_21_ ( .D(n740), .CK(clk), .RN(rstx), .Q(
        fu_ALU_o1reg[21]) );
  DFFRQX4 inst_decoder_rf_RF_rd_opc_reg_reg_0_ ( .D(n1181), .CK(clk), .RN(rstx), .Q(rf_RF_r1opcode_wire[0]) );
  DFFRQX4 inst_fetch_instruction_reg_reg_38_ ( .D(n1195), .CK(clk), .RN(rstx), 
        .Q(inst_decoder_instructionword_wire[38]) );
  DFFRQX4 fu_LSU_o1shadow_reg_reg_0_ ( .D(n1132), .CK(clk), .RN(rstx), .Q(
        fu_LSU_o1shadow_reg_0_) );
  DFFRQX4 fu_LSU_o1shadow_reg_reg_1_ ( .D(n1032), .CK(clk), .RN(rstx), .Q(
        fu_LSU_o1shadow_reg_1_) );
  DFFRQX4 inst_decoder_rf_BOOL_rd_opc_reg_reg_0_ ( .D(n1185), .CK(clk), .RN(
        rstx), .Q(rf_BOOL_r1opcode_wire_0_) );
  DFFRQX4 inst_decoder_fu_gcu_pc_load_reg_reg ( .D(n1135), .CK(clk), .RN(rstx), 
        .Q(inst_fetch_pc_load_wire) );
  INVX2 U1146 ( .A(inst_decoder_instructionword_wire[39]), .Y(n603) );
  INVX2 U1273 ( .A(rf_RF_r1opcode_wire[1]), .Y(n582) );
  INVX2 fu_ALU_fu_arch_U389 ( .A(fu_ALU_o1reg[16]), .Y(fu_ALU_fu_arch_n617) );
  NAND2X2 U1275 ( .A(ic_socket_RF_o1_bus_cntrl_wire_0_), .B(
        rf_RF_r1opcode_wire[1]), .Y(n631) );
  INVX2 U1017 ( .A(rf_RF_t1opcode_wire[2]), .Y(n548) );
  INVX2 U1141 ( .A(rf_BOOL_reg_0__0_), .Y(n602) );
  NAND2X2 U1016 ( .A(inst_decoder_N232), .B(inst_decoder_N230), .Y(n542) );
  INVX2 U1123 ( .A(inst_decoder_instructionword_wire[36]), .Y(n573) );
  NOR2X2 U911 ( .A(busy), .B(inst_fetch_pc_load_wire), .Y(n275) );
  NOR2X2 U876 ( .A(n458), .B(n459), .Y(n496) );
  NAND2X2 U877 ( .A(fu_LSU_status_addr_reg_1__3_), .B(n459), .Y(n493) );
  AO22X2 U701 ( .A0(n2258), .A1(ic_simm_B1_wire[2]), .B0(n2256), .B1(
        ic_socket_LIFTING_o1_data0_wire[2]), .Y(n402) );
  AO22X2 U672 ( .A0(n2258), .A1(ic_simm_B1_wire[3]), .B0(n2256), .B1(
        ic_socket_LIFTING_o1_data0_wire[3]), .Y(n392) );
  AO22X2 U479 ( .A0(n2258), .A1(ic_simm_B1_wire[10]), .B0(n2256), .B1(
        ic_socket_LIFTING_o1_data0_wire[10]), .Y(n315) );
  AO22X2 U450 ( .A0(n2258), .A1(ic_simm_B1_wire[11]), .B0(n2256), .B1(
        ic_socket_LIFTING_o1_data0_wire[11]), .Y(n304) );
  AO22X2 U537 ( .A0(n2258), .A1(ic_simm_B1_wire[8]), .B0(n2256), .B1(
        ic_socket_LIFTING_o1_data0_wire[8]), .Y(n341) );
  AO22X2 U645 ( .A0(n2258), .A1(ic_simm_B1_wire[4]), .B0(n2256), .B1(
        ic_socket_LIFTING_o1_data0_wire[4]), .Y(n382) );
  AO22X2 U1159 ( .A0(n2256), .A1(ic_socket_LIFTING_o1_data0_wire[0]), .B0(
        n2187), .B1(ic_socket_lsu_o1_data0_wire[0]), .Y(n613) );
  AO22X2 U421 ( .A0(n2258), .A1(ic_simm_B1_wire[12]), .B0(n2256), .B1(
        ic_socket_LIFTING_o1_data0_wire[12]), .Y(n293) );
  AO22X2 U564 ( .A0(n2258), .A1(ic_simm_B1_wire[7]), .B0(n2256), .B1(
        ic_socket_LIFTING_o1_data0_wire[7]), .Y(n352) );
  AO22X2 U618 ( .A0(n2258), .A1(ic_simm_B1_wire[5]), .B0(n2256), .B1(
        ic_socket_LIFTING_o1_data0_wire[5]), .Y(n372) );
  AO22X2 U591 ( .A0(n2258), .A1(ic_simm_B1_wire[6]), .B0(n2256), .B1(
        ic_socket_LIFTING_o1_data0_wire[6]), .Y(n362) );
  AO22X2 U508 ( .A0(n2258), .A1(ic_simm_B1_wire[9]), .B0(n2256), .B1(
        ic_socket_LIFTING_o1_data0_wire[9]), .Y(n328) );
  AO22X2 U392 ( .A0(n2258), .A1(ic_simm_B1_wire[13]), .B0(n2256), .B1(
        ic_socket_LIFTING_o1_data0_wire[13]), .Y(n282) );
  AOI222X2 U47 ( .A0(ic_socket_lsu_o1_data0_wire[29]), .A1(n2187), .B0(n59), 
        .B1(rf_RF_reg_2__29_), .C0(n2256), .C1(
        ic_socket_LIFTING_o1_data0_wire[29]), .Y(n71) );
  AOI222X2 U68 ( .A0(ic_socket_lsu_o1_data0_wire[28]), .A1(n2187), .B0(n59), 
        .B1(rf_RF_reg_2__28_), .C0(n2256), .C1(
        ic_socket_LIFTING_o1_data0_wire[28]), .Y(n83) );
  AO22X2 U929 ( .A0(n2258), .A1(ic_simm_B1_wire[14]), .B0(n2256), .B1(
        ic_socket_LIFTING_o1_data0_wire[14]), .Y(n511) );
  AOI222X2 U26 ( .A0(ic_socket_lsu_o1_data0_wire[30]), .A1(n2187), .B0(n59), 
        .B1(rf_RF_reg_2__30_), .C0(n2256), .C1(
        ic_socket_LIFTING_o1_data0_wire[30]), .Y(n55) );
  INVX6 fu_ALU_fu_arch_U687 ( .A(n2176), .Y(fu_ALU_fu_arch_n335) );
  INVX2 U1140 ( .A(n601), .Y(n559) );
  AOI22X2 U905 ( .A0(busy), .A1(inst_fetch_pc_reg_0_), .B0(n2114), .B1(
        inst_fetch_increased_pc_0_), .Y(n505) );
  AOI22X2 U682 ( .A0(busy), .A1(inst_fetch_pc_reg_2_), .B0(n2114), .B1(
        inst_fetch_increased_pc_2_), .Y(n396) );
  AO22X2 U1282 ( .A0(n2258), .A1(ic_simm_B1_wire[1]), .B0(n2256), .B1(
        ic_socket_LIFTING_o1_data0_wire[1]), .Y(n632) );
  AOI22X2 U746 ( .A0(busy), .A1(inst_fetch_pc_reg_1_), .B0(n2114), .B1(
        inst_fetch_increased_pc_1_), .Y(n410) );
  AOI2BB2X2 U900 ( .B0(inst_fetch_ra_load_wire), .B1(n2208), .A0N(n1282), 
        .A1N(inst_fetch_pc_opcode_wire_0_), .Y(n266) );
  AOI22X2 U504 ( .A0(ic_socket_lsu_o1_bus_cntrl_wire_0_), .A1(
        ic_socket_lsu_o1_data0_wire[9]), .B0(n2221), .B1(rf_RF_reg_4__9_), .Y(
        n327) );
  AOI22X2 U475 ( .A0(ic_socket_lsu_o1_bus_cntrl_wire_0_), .A1(
        ic_socket_lsu_o1_data0_wire[10]), .B0(n2221), .B1(rf_RF_reg_4__10_), 
        .Y(n314) );
  AOI22X2 U446 ( .A0(n2187), .A1(ic_socket_lsu_o1_data0_wire[11]), .B0(n2221), 
        .B1(rf_RF_reg_4__11_), .Y(n303) );
  NAND2X2 fu_ALU_fu_arch_U678 ( .A(n1768), .B(fu_ALU_fu_arch_n335), .Y(
        fu_ALU_fu_arch_n379) );
  AOI22X2 U653 ( .A0(busy), .A1(inst_fetch_pc_reg_3_), .B0(n2114), .B1(
        inst_fetch_increased_pc_3_), .Y(n386) );
  INVX2 U818 ( .A(n470), .Y(n456) );
  NAND2X2 U760 ( .A(n132), .B(n115), .Y(n319) );
  AOI22X2 U587 ( .A0(ic_socket_lsu_o1_bus_cntrl_wire_0_), .A1(
        ic_socket_lsu_o1_data0_wire[6]), .B0(n2221), .B1(rf_RF_reg_4__6_), .Y(
        n361) );
  AOI22X2 U668 ( .A0(n2187), .A1(ic_socket_lsu_o1_data0_wire[3]), .B0(n2221), 
        .B1(rf_RF_reg_4__3_), .Y(n391) );
  AOI22X2 U925 ( .A0(n2187), .A1(ic_socket_lsu_o1_data0_wire[14]), .B0(n2221), 
        .B1(rf_RF_reg_4__14_), .Y(n510) );
  AOI22X2 U560 ( .A0(ic_socket_lsu_o1_bus_cntrl_wire_0_), .A1(
        ic_socket_lsu_o1_data0_wire[7]), .B0(n2221), .B1(rf_RF_reg_4__7_), .Y(
        n351) );
  NAND2X2 fu_ALU_fu_arch_U552 ( .A(fu_ALU_fu_arch_n723), .B(n2167), .Y(
        fu_ALU_fu_arch_n633) );
  AOI22X2 U697 ( .A0(n2187), .A1(ic_socket_lsu_o1_data0_wire[2]), .B0(n2221), 
        .B1(rf_RF_reg_4__2_), .Y(n401) );
  AOI22X2 U614 ( .A0(n2187), .A1(ic_socket_lsu_o1_data0_wire[5]), .B0(n2221), 
        .B1(rf_RF_reg_4__5_), .Y(n371) );
  AOI22X2 U533 ( .A0(n2187), .A1(ic_socket_lsu_o1_data0_wire[8]), .B0(n2221), 
        .B1(rf_RF_reg_4__8_), .Y(n340) );
  AOI22X2 U641 ( .A0(n2187), .A1(ic_socket_lsu_o1_data0_wire[4]), .B0(n2221), 
        .B1(rf_RF_reg_4__4_), .Y(n381) );
  NAND2X2 U141 ( .A(fu_LSU_o1shadow_reg_0_), .B(n132), .Y(n125) );
  AOI22X2 U535 ( .A0(n2219), .A1(rf_RF_reg_0__8_), .B0(n2216), .B1(
        rf_RF_reg_1__8_), .Y(n338) );
  AOI22X2 U562 ( .A0(n2220), .A1(rf_RF_reg_0__7_), .B0(n2216), .B1(
        rf_RF_reg_1__7_), .Y(n349) );
  AOI22X2 U286 ( .A0(n2214), .A1(rf_RF_reg_2__18_), .B0(n2256), .B1(
        ic_socket_LIFTING_o1_data0_wire[18]), .Y(n213) );
  AOI22X2 U699 ( .A0(n2220), .A1(rf_RF_reg_0__2_), .B0(n2215), .B1(
        rf_RF_reg_1__2_), .Y(n399) );
  AOI22X2 U333 ( .A0(n2214), .A1(rf_RF_reg_2__16_), .B0(n2256), .B1(
        ic_socket_LIFTING_o1_data0_wire[16]), .Y(n246) );
  AOI22X2 U308 ( .A0(n2214), .A1(rf_RF_reg_2__17_), .B0(n2256), .B1(
        ic_socket_LIFTING_o1_data0_wire[17]), .Y(n226) );
  AOI22X2 U355 ( .A0(n2214), .A1(rf_RF_reg_2__15_), .B0(n2256), .B1(
        ic_socket_LIFTING_o1_data0_wire[15]), .Y(n258) );
  AOI22X2 U477 ( .A0(n2220), .A1(rf_RF_reg_0__10_), .B0(n2216), .B1(
        rf_RF_reg_1__10_), .Y(n312) );
  AOI22X2 U222 ( .A0(n2214), .A1(rf_RF_reg_2__21_), .B0(n2256), .B1(
        ic_socket_LIFTING_o1_data0_wire[21]), .Y(n175) );
  AOI222X2 U133 ( .A0(ic_socket_lsu_o1_data0_wire[25]), .A1(
        ic_socket_lsu_o1_bus_cntrl_wire_0_), .B0(n2214), .B1(rf_RF_reg_2__25_), 
        .C0(n2256), .C1(ic_socket_LIFTING_o1_data0_wire[25]), .Y(n121) );
  OAI21X4 fu_ALU_fu_arch_U399 ( .A0(fu_ALU_fu_arch_n631), .A1(n1767), .B0(
        fu_ALU_fu_arch_n633), .Y(fu_ALU_fu_arch_n290) );
  AOI22X2 U417 ( .A0(ic_socket_lsu_o1_bus_cntrl_wire_0_), .A1(
        ic_socket_lsu_o1_data0_wire[12]), .B0(n2222), .B1(rf_RF_reg_4__12_), 
        .Y(n292) );
  NAND2X2 fu_ALU_fu_arch_U625 ( .A(n2201), .B(n2161), .Y(fu_ALU_fu_arch_n687)
         );
  AOI22X2 U419 ( .A0(n2219), .A1(rf_RF_reg_0__12_), .B0(n2216), .B1(
        rf_RF_reg_1__12_), .Y(n290) );
  NAND2X2 fu_ALU_fu_arch_U558 ( .A(n2201), .B(fu_ALU_fu_arch_sub_200_B_8_), 
        .Y(fu_ALU_fu_arch_n327) );
  NAND2X2 fu_ALU_fu_arch_U665 ( .A(n2201), .B(n2132), .Y(fu_ALU_fu_arch_n370)
         );
  AOI22X2 U616 ( .A0(n2220), .A1(rf_RF_reg_0__5_), .B0(n2216), .B1(
        rf_RF_reg_1__5_), .Y(n369) );
  AOI22X2 U1268 ( .A0(n2187), .A1(ic_socket_lsu_o1_data0_wire[1]), .B0(n2222), 
        .B1(rf_RF_reg_4__1_), .Y(n630) );
  AOI22X2 U1276 ( .A0(n2220), .A1(rf_RF_reg_0__1_), .B0(n2215), .B1(
        rf_RF_reg_1__1_), .Y(n628) );
  NAND2X2 fu_ALU_fu_arch_U444 ( .A(n2201), .B(fu_ALU_fu_arch_sub_200_B_11_), 
        .Y(fu_ALU_fu_arch_n546) );
  NAND2X2 fu_ALU_fu_arch_U640 ( .A(n2201), .B(fu_ALU_o1reg[6]), .Y(
        fu_ALU_fu_arch_n689) );
  INVX6 fu_ALU_fu_arch_U551 ( .A(fu_ALU_fu_arch_n633), .Y(fu_ALU_fu_arch_n128)
         );
  NAND2X2 fu_ALU_fu_arch_U471 ( .A(n2201), .B(n2153), .Y(fu_ALU_fu_arch_n605)
         );
  NAND2X2 fu_ALU_fu_arch_U451 ( .A(n2201), .B(fu_ALU_o1reg[3]), .Y(
        fu_ALU_fu_arch_n550) );
  AOI222X2 U159 ( .A0(ic_socket_lsu_o1_data0_wire[24]), .A1(
        ic_socket_lsu_o1_bus_cntrl_wire_0_), .B0(n2214), .B1(rf_RF_reg_2__24_), 
        .C0(n2256), .C1(ic_socket_LIFTING_o1_data0_wire[24]), .Y(n137) );
  AOI22X2 U506 ( .A0(n2219), .A1(rf_RF_reg_0__9_), .B0(n2216), .B1(
        rf_RF_reg_1__9_), .Y(n325) );
  AOI22X2 U243 ( .A0(n2214), .A1(rf_RF_reg_2__20_), .B0(n2256), .B1(
        ic_socket_LIFTING_o1_data0_wire[20]), .Y(n187) );
  CLKNAND2X2 fu_ALU_fu_arch_U309 ( .A(n2201), .B(n2166), .Y(
        fu_ALU_fu_arch_n553) );
  AOI22X2 U626 ( .A0(busy), .A1(inst_fetch_pc_reg_4_), .B0(n2114), .B1(
        inst_fetch_increased_pc_4_), .Y(n376) );
  AOI22X2 U201 ( .A0(n2214), .A1(rf_RF_reg_2__22_), .B0(n2256), .B1(
        ic_socket_LIFTING_o1_data0_wire[22]), .Y(n163) );
  NAND2X2 fu_ALU_fu_arch_U682 ( .A(n2201), .B(fu_ALU_fu_arch_sub_200_B_18_), 
        .Y(fu_ALU_fu_arch_n524) );
  NAND2X2 fu_ALU_fu_arch_U464 ( .A(n2201), .B(n2138), .Y(fu_ALU_fu_arch_n422)
         );
  AOI22X2 U388 ( .A0(n2187), .A1(ic_socket_lsu_o1_data0_wire[13]), .B0(n2222), 
        .B1(rf_RF_reg_4__13_), .Y(n281) );
  NAND2X2 fu_ALU_fu_arch_U630 ( .A(n2201), .B(fu_ALU_fu_arch_sub_200_B_14_), 
        .Y(fu_ALU_fu_arch_n623) );
  AOI22X2 U390 ( .A0(n2219), .A1(rf_RF_reg_0__13_), .B0(n2216), .B1(
        rf_RF_reg_1__13_), .Y(n279) );
  AOI22X2 U264 ( .A0(n2214), .A1(rf_RF_reg_2__19_), .B0(
        ic_socket_LIFTING_o1_bus_cntrl_wire_0_), .B1(
        ic_socket_LIFTING_o1_data0_wire[19]), .Y(n199) );
  AOI22X2 U180 ( .A0(n2214), .A1(rf_RF_reg_2__23_), .B0(n2256), .B1(
        ic_socket_LIFTING_o1_data0_wire[23]), .Y(n151) );
  NAND2X2 fu_ALU_fu_arch_U458 ( .A(n2201), .B(fu_ALU_fu_arch_sub_200_B_19_), 
        .Y(fu_ALU_fu_arch_n517) );
  NAND2X2 fu_ALU_fu_arch_U434 ( .A(n2201), .B(fu_ALU_fu_arch_sub_200_B_27_), 
        .Y(fu_ALU_fu_arch_n350) );
  NAND2X2 fu_ALU_fu_arch_U699 ( .A(n2201), .B(fu_ALU_fu_arch_sub_200_B_22_), 
        .Y(fu_ALU_fu_arch_n446) );
  AOI22X2 U307 ( .A0(n2217), .A1(rf_RF_reg_3__17_), .B0(n2216), .B1(
        rf_RF_reg_1__17_), .Y(n227) );
  NOR2X2 fu_ALU_fu_arch_U703 ( .A(fu_ALU_fu_arch_n274), .B(n1851), .Y(
        fu_ALU_fu_arch_n737) );
  AOI22X2 U263 ( .A0(n2217), .A1(rf_RF_reg_3__19_), .B0(n2215), .B1(
        rf_RF_reg_1__19_), .Y(n200) );
  AOI22X2 U132 ( .A0(n2217), .A1(rf_RF_reg_3__25_), .B0(n2215), .B1(
        rf_RF_reg_1__25_), .Y(n122) );
  AOI22X2 U67 ( .A0(n2217), .A1(rf_RF_reg_3__28_), .B0(n2215), .B1(
        rf_RF_reg_1__28_), .Y(n84) );
  AOI22X2 U332 ( .A0(n2217), .A1(rf_RF_reg_3__16_), .B0(n2216), .B1(
        rf_RF_reg_1__16_), .Y(n247) );
  AOI22X2 U389 ( .A0(n2214), .A1(rf_RF_reg_2__13_), .B0(n2217), .B1(
        rf_RF_reg_3__13_), .Y(n280) );
  AOI22X2 U179 ( .A0(n2217), .A1(rf_RF_reg_3__23_), .B0(n2215), .B1(
        rf_RF_reg_1__23_), .Y(n152) );
  AOI22X2 U221 ( .A0(n2217), .A1(rf_RF_reg_3__21_), .B0(n2215), .B1(
        rf_RF_reg_1__21_), .Y(n176) );
  AOI22X2 U158 ( .A0(n2217), .A1(rf_RF_reg_3__24_), .B0(n2215), .B1(
        rf_RF_reg_1__24_), .Y(n138) );
  AOI22X2 U200 ( .A0(n2217), .A1(rf_RF_reg_3__22_), .B0(n2215), .B1(
        rf_RF_reg_1__22_), .Y(n164) );
  NOR2X2 fu_ALU_fu_arch_U378 ( .A(n2203), .B(fu_ALU_fu_arch_n108), .Y(
        fu_ALU_fu_arch_n391) );
  AOI22X2 U599 ( .A0(busy), .A1(inst_fetch_pc_reg_5_), .B0(n2114), .B1(
        inst_fetch_increased_pc_5_), .Y(n366) );
  NOR2X2 U899 ( .A(inst_fetch_ra_load_wire), .B(n2115), .Y(n267) );
  INVX2 fu_ALU_fu_arch_U578 ( .A(fu_ALU_fu_arch_n592), .Y(fu_ALU_fu_arch_n499)
         );
  CLKNAND2X2 fu_ALU_fu_arch_U588 ( .A(n2197), .B(fu_ALU_fu_arch_sub_200_B_18_), 
        .Y(fu_ALU_fu_arch_n733) );
  NOR2X2 fu_ALU_fu_arch_U417 ( .A(n2179), .B(n2195), .Y(fu_ALU_fu_arch_n647)
         );
  AOI22X2 U572 ( .A0(busy), .A1(inst_fetch_pc_reg_6_), .B0(n2114), .B1(
        inst_fetch_increased_pc_6_), .Y(n356) );
  AOI22X2 fu_ALU_fu_arch_U429 ( .A0(n2198), .A1(fu_ALU_o1reg[14]), .B0(n2201), 
        .B1(n2157), .Y(fu_ALU_fu_arch_n654) );
  NAND2X2 fu_ALU_fu_arch_U561 ( .A(n2197), .B(fu_ALU_o1reg[6]), .Y(
        fu_ALU_fu_arch_n326) );
  NAND2X2 fu_ALU_fu_arch_U574 ( .A(n2197), .B(n2132), .Y(fu_ALU_fu_arch_n729)
         );
  NAND2X2 fu_ALU_fu_arch_U463 ( .A(n2197), .B(fu_ALU_fu_arch_sub_200_B_21_), 
        .Y(fu_ALU_fu_arch_n670) );
  CLKNAND2X2 fu_ALU_fu_arch_U594 ( .A(n2197), .B(fu_ALU_o1reg[10]), .Y(
        fu_ALU_fu_arch_n735) );
  NOR2X2 fu_ALU_fu_arch_U201 ( .A(n2135), .B(n2195), .Y(fu_ALU_fu_arch_n429)
         );
  NAND2X2 U24 ( .A(n55), .B(n56), .Y(n54) );
  OAI211X2 U331 ( .A0(n149), .A1(n245), .B0(n246), .C0(n247), .Y(n244) );
  AOI22X2 fu_ALU_fu_arch_U349 ( .A0(n2198), .A1(fu_ALU_fu_arch_sub_200_B_18_), 
        .B0(n2201), .B1(fu_ALU_o1reg[16]), .Y(fu_ALU_fu_arch_n588) );
  NOR2X2 fu_ALU_fu_arch_U291 ( .A(fu_ALU_o1reg[20]), .B(n2195), .Y(
        fu_ALU_fu_arch_n532) );
  NAND2X2 U157 ( .A(n137), .B(n138), .Y(n136) );
  OAI211X2 U199 ( .A0(n149), .A1(n162), .B0(n163), .C0(n164), .Y(n161) );
  NAND2X2 U87 ( .A(n95), .B(n96), .Y(n94) );
  NOR2X2 fu_ALU_fu_arch_U272 ( .A(fu_ALU_fu_arch_sub_200_B_21_), .B(n2195), 
        .Y(fu_ALU_fu_arch_n514) );
  OAI211X2 U306 ( .A0(n149), .A1(n225), .B0(n226), .C0(n227), .Y(n224) );
  NOR2X2 fu_ALU_fu_arch_U204 ( .A(fu_ALU_o1reg[25]), .B(n2196), .Y(
        fu_ALU_fu_arch_n433) );
  NOR2X2 fu_ALU_fu_arch_U253 ( .A(n2141), .B(n2195), .Y(fu_ALU_fu_arch_n494)
         );
  NOR2X2 fu_ALU_fu_arch_U115 ( .A(fu_ALU_fu_arch_sub_200_B_30_), .B(n2196), 
        .Y(fu_ALU_fu_arch_n301) );
  OAI211X2 U284 ( .A0(n149), .A1(n212), .B0(n213), .C0(n214), .Y(n211) );
  NAND2X2 U109 ( .A(n108), .B(n109), .Y(n107) );
  OAI211X2 U241 ( .A0(n149), .A1(n186), .B0(n187), .C0(n188), .Y(n185) );
  NAND2X2 U45 ( .A(n71), .B(n72), .Y(n70) );
  NAND2X2 fu_ALU_fu_arch_U379 ( .A(n2105), .B(fu_ALU_fu_arch_n612), .Y(
        fu_ALU_fu_arch_n601) );
  OAI211X2 U942 ( .A0(n149), .A1(n491), .B0(n517), .C0(n518), .Y(n516) );
  NAND2X4 fu_ALU_fu_arch_U165 ( .A(fu_ALU_fu_arch_n278), .B(n1851), .Y(
        fu_ALU_fu_arch_n270) );
  NAND2X2 U131 ( .A(n121), .B(n122), .Y(n120) );
  OAI2B11X2 U353 ( .A1N(ic_socket_lsu_o1_data0_wire[15]), .A0(n149), .B0(n258), 
        .C0(n259), .Y(n257) );
  NAND2X2 fu_ALU_fu_arch_U697 ( .A(n2197), .B(n2144), .Y(fu_ALU_fu_arch_n767)
         );
  OAI211X2 U220 ( .A0(n149), .A1(n174), .B0(n175), .C0(n176), .Y(n173) );
  NAND2X2 fu_ALU_fu_arch_U516 ( .A(n2197), .B(n2166), .Y(fu_ALU_fu_arch_n259)
         );
  NAND2X4 fu_ALU_fu_arch_U637 ( .A(n2197), .B(n2181), .Y(fu_ALU_fu_arch_n619)
         );
  OAI211X2 U262 ( .A0(n149), .A1(n198), .B0(n199), .C0(n200), .Y(n197) );
  NAND2X2 U66 ( .A(n83), .B(n84), .Y(n82) );
  OAI211X2 U178 ( .A0(n149), .A1(n150), .B0(n151), .C0(n152), .Y(n148) );
  AOI22X2 fu_ALU_fu_arch_U247 ( .A0(fu_ALU_fu_arch_n284), .A1(fu_ALU_o1reg[19]), .B0(n2201), .B1(n2144), .Y(fu_ALU_fu_arch_n486) );
  AOI211X4 fu_ALU_fu_arch_U339 ( .A0(n2188), .A1(n2149), .B0(
        fu_ALU_fu_arch_n583), .C0(n2190), .Y(fu_ALU_fu_arch_n581) );
  AOI22X2 fu_ALU_fu_arch_U514 ( .A0(n2198), .A1(fu_ALU_o1reg[11]), .B0(n2202), 
        .B1(fu_ALU_fu_arch_sub_200_B_8_), .Y(fu_ALU_fu_arch_n702) );
  NAND2X2 fu_ALU_fu_arch_U690 ( .A(n2200), .B(fu_ALU_o1reg[21]), .Y(
        fu_ALU_fu_arch_n487) );
  AOI22X2 fu_ALU_fu_arch_U559 ( .A0(n2198), .A1(n2161), .B0(n2202), .B1(n2166), 
        .Y(fu_ALU_fu_arch_n724) );
  AOI22X2 fu_ALU_fu_arch_U495 ( .A0(n2198), .A1(fu_ALU_o1reg[12]), .B0(n2200), 
        .B1(fu_ALU_o1reg[11]), .Y(fu_ALU_fu_arch_n686) );
  AOI32X2 fu_ALU_fu_arch_U326 ( .A0(n2147), .A1(n2146), .A2(n1762), .B0(n2190), 
        .B1(n2147), .Y(fu_ALU_fu_arch_n569) );
  NAND2X2 fu_ALU_fu_arch_U629 ( .A(n2202), .B(n2153), .Y(fu_ALU_fu_arch_n589)
         );
  NAND2X2 fu_ALU_fu_arch_U624 ( .A(n2202), .B(fu_ALU_fu_arch_sub_200_B_11_), 
        .Y(fu_ALU_fu_arch_n655) );
  AOI22X2 fu_ALU_fu_arch_U497 ( .A0(n2198), .A1(fu_ALU_fu_arch_sub_200_B_8_), 
        .B0(n2200), .B1(n2166), .Y(fu_ALU_fu_arch_n688) );
  NAND2X2 fu_ALU_fu_arch_U694 ( .A(n2202), .B(n2138), .Y(fu_ALU_fu_arch_n412)
         );
  AOI22X2 fu_ALU_fu_arch_U524 ( .A0(n2198), .A1(fu_ALU_fu_arch_sub_200_B_11_), 
        .B0(n2202), .B1(fu_ALU_fu_arch_sub_200_B_14_), .Y(fu_ALU_fu_arch_n705)
         );
  INVX2 fu_ALU_fu_arch_U636 ( .A(fu_ALU_fu_arch_n619), .Y(fu_ALU_fu_arch_n459)
         );
  AOI22X2 fu_ALU_fu_arch_U452 ( .A0(n2198), .A1(fu_ALU_fu_arch_sub_200_B_5_), 
        .B0(n2200), .B1(fu_ALU_fu_arch_sub_200_B_4_), .Y(fu_ALU_fu_arch_n668)
         );
  NOR2X2 fu_ALU_fu_arch_U381 ( .A(fu_ALU_fu_arch_n468), .B(fu_ALU_fu_arch_n108), .Y(fu_ALU_fu_arch_n394) );
  AOI22X2 U545 ( .A0(busy), .A1(inst_fetch_pc_reg_7_), .B0(n2114), .B1(
        inst_fetch_increased_pc_7_), .Y(n346) );
  AOI22X2 fu_ALU_fu_arch_U562 ( .A0(n2095), .A1(fu_ALU_fu_arch_sub_200_B_4_), 
        .B0(n2200), .B1(fu_ALU_fu_arch_sub_200_B_5_), .Y(fu_ALU_fu_arch_n725)
         );
  INVX2 U951 ( .A(n523), .Y(n1099) );
  INVX2 fu_ALU_fu_arch_U533 ( .A(fu_ALU_fu_arch_n283), .Y(fu_ALU_fu_arch_n635)
         );
  AOI32X2 fu_ALU_fu_arch_U364 ( .A0(n2150), .A1(fu_ALU_fu_arch_n522), .A2(
        n1762), .B0(n2190), .B1(n2150), .Y(fu_ALU_fu_arch_n602) );
  NAND2X2 fu_ALU_fu_arch_U531 ( .A(n2200), .B(fu_ALU_fu_arch_lt_gt_188_A_28_), 
        .Y(fu_ALU_fu_arch_n708) );
  NAND2X2 fu_ALU_fu_arch_U513 ( .A(n2200), .B(fu_ALU_o1reg[10]), .Y(
        fu_ALU_fu_arch_n547) );
  OAI211X2 fu_ALU_fu_arch_U563 ( .A0(n2162), .A1(n2196), .B0(
        fu_ALU_fu_arch_n726), .C0(n2092), .Y(fu_ALU_fu_arch_n719) );
  AOI22X2 fu_ALU_fu_arch_U330 ( .A0(n2197), .A1(fu_ALU_fu_arch_sub_200_B_19_), 
        .B0(n2202), .B1(fu_ALU_o1reg[16]), .Y(fu_ALU_fu_arch_n571) );
  NAND2X2 fu_ALU_fu_arch_U461 ( .A(n2200), .B(fu_ALU_o1reg[22]), .Y(
        fu_ALU_fu_arch_n467) );
  AOI211X4 fu_ALU_fu_arch_U416 ( .A0(n2188), .A1(n2179), .B0(
        fu_ALU_fu_arch_n647), .C0(n2190), .Y(fu_ALU_fu_arch_n645) );
  AOI22X2 fu_ALU_fu_arch_U585 ( .A0(n2201), .A1(n2151), .B0(n2200), .B1(n2153), 
        .Y(fu_ALU_fu_arch_n730) );
  OAI211X2 fu_ALU_fu_arch_U100 ( .A0(n2199), .A1(fu_ALU_fu_arch_n270), .B0(
        fu_ALU_fu_arch_n271), .C0(n2092), .Y(fu_ALU_fu_arch_n268) );
  INVX2 fu_ALU_fu_arch_U39 ( .A(fu_ALU_fu_arch_n153), .Y(fu_ALU_fu_arch_n125)
         );
  NAND2X2 fu_ALU_fu_arch_U540 ( .A(n2200), .B(n2144), .Y(fu_ALU_fu_arch_n712)
         );
  AOI22X2 fu_ALU_fu_arch_U445 ( .A0(n2202), .A1(fu_ALU_o1reg[10]), .B0(n2200), 
        .B1(fu_ALU_o1reg[12]), .Y(fu_ALU_fu_arch_n666) );
  AOI22X2 fu_ALU_fu_arch_U683 ( .A0(n2197), .A1(n2151), .B0(n2202), .B1(
        fu_ALU_fu_arch_sub_200_B_19_), .Y(fu_ALU_fu_arch_n766) );
  NAND2X2 fu_ALU_fu_arch_U447 ( .A(n2202), .B(n2168), .Y(fu_ALU_fu_arch_n253)
         );
  AOI22X2 fu_ALU_fu_arch_U510 ( .A0(n2198), .A1(n2173), .B0(n2181), .B1(n2202), 
        .Y(fu_ALU_fu_arch_n701) );
  NAND2X2 fu_ALU_fu_arch_U462 ( .A(n2202), .B(fu_ALU_o1reg[24]), .Y(
        fu_ALU_fu_arch_n393) );
  AOI22X2 fu_ALU_fu_arch_U448 ( .A0(n2201), .A1(n2166), .B0(n2200), .B1(
        fu_ALU_o1reg[8]), .Y(fu_ALU_fu_arch_n667) );
  NAND2X2 fu_ALU_fu_arch_U457 ( .A(n2200), .B(fu_ALU_fu_arch_sub_200_B_18_), 
        .Y(fu_ALU_fu_arch_n572) );
  AOI211X4 fu_ALU_fu_arch_U319 ( .A0(n2188), .A1(n2147), .B0(
        fu_ALU_fu_arch_n566), .C0(n2190), .Y(fu_ALU_fu_arch_n564) );
  AOI22X2 fu_ALU_fu_arch_U230 ( .A0(n2197), .A1(fu_ALU_o1reg[23]), .B0(n2202), 
        .B1(n2144), .Y(fu_ALU_fu_arch_n466) );
  AOI211X4 fu_ALU_fu_arch_U466 ( .A0(n2156), .A1(n2188), .B0(n2190), .C0(
        fu_ALU_fu_arch_n672), .Y(fu_ALU_fu_arch_n671) );
  NAND2X2 fu_ALU_fu_arch_U543 ( .A(n2200), .B(n2136), .Y(fu_ALU_fu_arch_n714)
         );
  AOI22X2 fu_ALU_fu_arch_U517 ( .A0(n2202), .A1(fu_ALU_o1reg[4]), .B0(n2200), 
        .B1(fu_ALU_o1reg[6]), .Y(fu_ALU_fu_arch_n703) );
  NAND2X2 fu_ALU_fu_arch_U509 ( .A(fu_ALU_fu_arch_sub_200_B_2_), .B(n2200), 
        .Y(fu_ALU_fu_arch_n551) );
  AOI22X2 fu_ALU_fu_arch_U589 ( .A0(n2201), .A1(fu_ALU_o1reg[20]), .B0(n2200), 
        .B1(fu_ALU_fu_arch_sub_200_B_19_), .Y(fu_ALU_fu_arch_n732) );
  AOI211X4 fu_ALU_fu_arch_U264 ( .A0(n2188), .A1(n2143), .B0(
        fu_ALU_fu_arch_n507), .C0(n2190), .Y(fu_ALU_fu_arch_n506) );
  AOI211X4 fu_ALU_fu_arch_U252 ( .A0(n2188), .A1(n2141), .B0(
        fu_ALU_fu_arch_n494), .C0(n2190), .Y(fu_ALU_fu_arch_n491) );
  AOI211X4 fu_ALU_fu_arch_U200 ( .A0(n2188), .A1(n2135), .B0(
        fu_ALU_fu_arch_n429), .C0(n2190), .Y(fu_ALU_fu_arch_n425) );
  AOI22X2 U611 ( .A0(ic_socket_gcu_o1_data0_wire[5]), .A1(n2115), .B0(n2116), 
        .B1(inst_fetch_increased_pc_5_), .Y(n367) );
  AOI22X2 U638 ( .A0(ic_socket_gcu_o1_data0_wire[4]), .A1(n2115), .B0(n2116), 
        .B1(inst_fetch_increased_pc_4_), .Y(n377) );
  AOI22X2 U895 ( .A0(ic_socket_gcu_o1_data0_wire[1]), .A1(n2115), .B0(n2116), 
        .B1(inst_fetch_increased_pc_1_), .Y(n502) );
  AOI22X2 U665 ( .A0(ic_socket_gcu_o1_data0_wire[3]), .A1(n2115), .B0(n2116), 
        .B1(inst_fetch_increased_pc_3_), .Y(n387) );
  AOI22X2 U694 ( .A0(ic_socket_gcu_o1_data0_wire[2]), .A1(n2115), .B0(n2116), 
        .B1(inst_fetch_increased_pc_2_), .Y(n397) );
  AOI22X2 U557 ( .A0(ic_socket_gcu_o1_data0_wire[7]), .A1(n2115), .B0(n2116), 
        .B1(inst_fetch_increased_pc_7_), .Y(n347) );
  AOI22X2 U584 ( .A0(ic_socket_gcu_o1_data0_wire[6]), .A1(n2115), .B0(n2116), 
        .B1(inst_fetch_increased_pc_6_), .Y(n357) );
  AOI22X2 fu_ALU_fu_arch_U277 ( .A0(n2202), .A1(fu_ALU_fu_arch_sub_200_B_18_), 
        .B0(n2200), .B1(n2144), .Y(fu_ALU_fu_arch_n516) );
  AOI22X2 fu_ALU_fu_arch_U213 ( .A0(n2197), .A1(n2136), .B0(n2200), .B1(
        fu_ALU_o1reg[23]), .Y(fu_ALU_fu_arch_n445) );
  AOI22X2 fu_ALU_fu_arch_U158 ( .A0(n2198), .A1(fu_ALU_o1reg[28]), .B0(n2200), 
        .B1(fu_ALU_fu_arch_sub_200_B_27_), .Y(fu_ALU_fu_arch_n369) );
  AOI22X2 U530 ( .A0(ic_socket_gcu_o1_data0_wire[8]), .A1(n2115), .B0(n2116), 
        .B1(inst_fetch_increased_pc_8_), .Y(n336) );
  AOI22X2 fu_ALU_fu_arch_U641 ( .A0(n2202), .A1(n2166), .B0(n2200), .B1(
        fu_ALU_fu_arch_sub_200_B_5_), .Y(fu_ALU_fu_arch_n758) );
  AOI22X2 fu_ALU_fu_arch_U283 ( .A0(n2197), .A1(n2144), .B0(n2200), .B1(
        fu_ALU_o1reg[19]), .Y(fu_ALU_fu_arch_n523) );
  NAND2X2 U975 ( .A(n2113), .B(n527), .Y(n534) );
  AOI22X2 U518 ( .A0(busy), .A1(inst_fetch_pc_reg_8_), .B0(n2114), .B1(
        inst_fetch_increased_pc_8_), .Y(n335) );
  AOI22X2 fu_ALU_fu_arch_U393 ( .A0(n2197), .A1(fu_ALU_o1reg[16]), .B0(n2200), 
        .B1(n2153), .Y(fu_ALU_fu_arch_n622) );
  AOI22X2 fu_ALU_fu_arch_U410 ( .A0(n2197), .A1(n2153), .B0(n2200), .B1(
        fu_ALU_o1reg[14]), .Y(fu_ALU_fu_arch_n639) );
  AOI22X2 fu_ALU_fu_arch_U367 ( .A0(n2202), .A1(fu_ALU_o1reg[14]), .B0(n2200), 
        .B1(n2151), .Y(fu_ALU_fu_arch_n604) );
  INVX2 U766 ( .A(n2113), .Y(n418) );
  AOI22X2 fu_ALU_fu_arch_U145 ( .A0(n2202), .A1(fu_ALU_o1reg[26]), .B0(n2200), 
        .B1(fu_ALU_o1reg[28]), .Y(fu_ALU_fu_arch_n348) );
  INVX2 fu_ALU_fu_arch_U688 ( .A(fu_ALU_fu_arch_n534), .Y(fu_ALU_fu_arch_n156)
         );
  AOI22X2 fu_ALU_fu_arch_U420 ( .A0(n2179), .A1(fu_ALU_fu_arch_n153), .B0(
        fu_ALU_fu_arch_n636), .B1(fu_ALU_fu_arch_n590), .Y(fu_ALU_fu_arch_n651) );
  INVX2 fu_ALU_fu_arch_U474 ( .A(fu_ALU_fu_arch_n434), .Y(fu_ALU_fu_arch_n337)
         );
  INVX2 U963 ( .A(n501), .Y(n500) );
  INVX2 fu_ALU_fu_arch_U275 ( .A(n1798), .Y(fu_ALU_fu_arch_n441) );
  AOI22X2 fu_ALU_fu_arch_U492 ( .A0(n1892), .A1(fu_ALU_fu_arch_n534), .B0(
        n1854), .B1(fu_ALU_fu_arch_n224), .Y(fu_ALU_fu_arch_n676) );
  AOI22X2 U489 ( .A0(busy), .A1(inst_fetch_pc_reg_9_), .B0(n2114), .B1(
        inst_fetch_increased_pc_9_), .Y(n322) );
  AOI22X2 U501 ( .A0(ic_socket_gcu_o1_data0_wire[9]), .A1(n2115), .B0(n2116), 
        .B1(inst_fetch_increased_pc_9_), .Y(n323) );
  AOI21X4 fu_ALU_fu_arch_U490 ( .A0(fu_ALU_fu_arch_n249), .A1(
        fu_ALU_fu_arch_n456), .B0(fu_ALU_fu_arch_n648), .Y(fu_ALU_fu_arch_n372) );
  AOI22X2 fu_ALU_fu_arch_U60 ( .A0(n1892), .A1(n1827), .B0(n1854), .B1(n1792), 
        .Y(fu_ALU_fu_arch_n181) );
  INVX2 fu_ALU_fu_arch_U347 ( .A(n1801), .Y(fu_ALU_fu_arch_n483) );
  AOI22X2 U460 ( .A0(busy), .A1(inst_fetch_pc_reg_10_), .B0(n2114), .B1(
        inst_fetch_increased_pc_10_), .Y(n309) );
  INVX2 fu_ALU_fu_arch_U321 ( .A(n1829), .Y(fu_ALU_fu_arch_n234) );
  AOI22X2 fu_ALU_fu_arch_U406 ( .A0(n2105), .A1(n1829), .B0(n2104), .B1(n1828), 
        .Y(fu_ALU_fu_arch_n638) );
  AOI22X2 fu_ALU_fu_arch_U582 ( .A0(n1892), .A1(n1831), .B0(n1854), .B1(n1827), 
        .Y(fu_ALU_fu_arch_n716) );
  AOI22X2 fu_ALU_fu_arch_U251 ( .A0(n2101), .A1(n1842), .B0(
        fu_ALU_fu_arch_n395), .B1(n1888), .Y(fu_ALU_fu_arch_n492) );
  AOI22X2 fu_ALU_fu_arch_U482 ( .A0(n2158), .A1(fu_ALU_fu_arch_n153), .B0(
        fu_ALU_fu_arch_n636), .B1(fu_ALU_fu_arch_n456), .Y(fu_ALU_fu_arch_n681) );
  NAND2X2 fu_ALU_fu_arch_U572 ( .A(fu_ALU_fu_arch_n249), .B(n1836), .Y(
        fu_ALU_fu_arch_n727) );
  AOI22X2 U472 ( .A0(ic_socket_gcu_o1_data0_wire[10]), .A1(n2115), .B0(n2116), 
        .B1(inst_fetch_increased_pc_10_), .Y(n310) );
  AOI22X2 fu_ALU_fu_arch_U411 ( .A0(n1833), .A1(n1834), .B0(n1854), .B1(n1839), 
        .Y(fu_ALU_fu_arch_n624) );
  AOI22X2 fu_ALU_fu_arch_U395 ( .A0(n2103), .A1(n1855), .B0(n1892), .B1(n1847), 
        .Y(fu_ALU_fu_arch_n626) );
  AOI22X2 fu_ALU_fu_arch_U171 ( .A0(n2100), .A1(n1793), .B0(
        fu_ALU_fu_arch_n333), .B1(fu_ALU_fu_arch_n285), .Y(fu_ALU_fu_arch_n390) );
  AOI22X2 fu_ALU_fu_arch_U430 ( .A0(n1833), .A1(n1827), .B0(n1854), .B1(n1831), 
        .Y(fu_ALU_fu_arch_n640) );
  OAI2BB2X2 fu_ALU_fu_arch_U263 ( .B0(fu_ALU_fu_arch_n506), .B1(n2142), .A0N(
        n1837), .A1N(fu_ALU_fu_arch_n395), .Y(fu_ALU_fu_arch_n505) );
  CLKINVX2 U764 ( .A(n206), .Y(n32) );
  AOI22X2 fu_ALU_fu_arch_U187 ( .A0(n2101), .A1(n1801), .B0(
        fu_ALU_fu_arch_n395), .B1(n1842), .Y(fu_ALU_fu_arch_n409) );
  AOI22X2 fu_ALU_fu_arch_U184 ( .A0(n2100), .A1(n1794), .B0(
        fu_ALU_fu_arch_n333), .B1(fu_ALU_fu_arch_n313), .Y(fu_ALU_fu_arch_n410) );
  AOI22X2 fu_ALU_fu_arch_U538 ( .A0(n2103), .A1(n1847), .B0(n1892), .B1(n1839), 
        .Y(fu_ALU_fu_arch_n692) );
  NAND2X2 fu_ALU_fu_arch_U293 ( .A(n1768), .B(fu_ALU_fu_arch_n533), .Y(
        fu_ALU_fu_arch_n228) );
  NOR2X2 U822 ( .A(n1806), .B(n2212), .Y(n474) );
  INVX2 fu_ALU_fu_arch_U328 ( .A(n1799), .Y(fu_ALU_fu_arch_n462) );
  OAI211X2 fu_ALU_fu_arch_U126 ( .A0(fu_ALU_fu_arch_n195), .A1(n2203), .B0(
        fu_ALU_fu_arch_n320), .C0(fu_ALU_fu_arch_n321), .Y(fu_ALU_fu_arch_n319) );
  OAI21X4 fu_ALU_fu_arch_U331 ( .A0(fu_ALU_fu_arch_n573), .A1(n1768), .B0(
        fu_ALU_fu_arch_n574), .Y(fu_ALU_fu_arch_n229) );
  AOI22X2 fu_ALU_fu_arch_U592 ( .A0(n2103), .A1(n1835), .B0(n1833), .B1(n1792), 
        .Y(fu_ALU_fu_arch_n715) );
  OAI21X4 fu_ALU_fu_arch_U231 ( .A0(fu_ALU_fu_arch_n468), .A1(
        fu_ALU_fu_arch_n283), .B0(fu_ALU_fu_arch_n469), .Y(fu_ALU_fu_arch_n179) );
  NAND2X2 fu_ALU_fu_arch_U242 ( .A(fu_ALU_fu_arch_n469), .B(
        fu_ALU_fu_arch_n437), .Y(fu_ALU_fu_arch_n177) );
  OAI211X2 fu_ALU_fu_arch_U250 ( .A0(fu_ALU_fu_arch_n491), .A1(n2140), .B0(
        fu_ALU_fu_arch_n492), .C0(n2102), .Y(fu_ALU_fu_arch_n490) );
  AOI22X2 U431 ( .A0(busy), .A1(inst_fetch_pc_reg_11_), .B0(n2114), .B1(
        inst_fetch_increased_pc_11_), .Y(n298) );
  AOI222X2 fu_ALU_fu_arch_U234 ( .A0(fu_ALU_o1reg[23]), .A1(
        fu_ALU_fu_arch_n473), .B0(n2101), .B1(n1841), .C0(fu_ALU_fu_arch_n395), 
        .C1(n1830), .Y(fu_ALU_fu_arch_n472) );
  AOI22X2 fu_ALU_fu_arch_U174 ( .A0(n2101), .A1(n1799), .B0(
        fu_ALU_fu_arch_n395), .B1(n1841), .Y(fu_ALU_fu_arch_n389) );
  AOI222X2 fu_ALU_fu_arch_U286 ( .A0(fu_ALU_o1reg[20]), .A1(
        fu_ALU_fu_arch_n528), .B0(n2100), .B1(n1840), .C0(fu_ALU_fu_arch_n395), 
        .C1(n1846), .Y(fu_ALU_fu_arch_n527) );
  OAI211X2 fu_ALU_fu_arch_U183 ( .A0(fu_ALU_fu_arch_n408), .A1(
        fu_ALU_fu_arch_n388), .B0(fu_ALU_fu_arch_n409), .C0(
        fu_ALU_fu_arch_n410), .Y(fu_ALU_fu_arch_n407) );
  AOI22X2 fu_ALU_fu_arch_U521 ( .A0(fu_ALU_fu_arch_n111), .A1(
        fu_ALU_fu_arch_n384), .B0(n1833), .B1(n1800), .Y(fu_ALU_fu_arch_n694)
         );
  INVX2 fu_ALU_fu_arch_U365 ( .A(n1796), .Y(fu_ALU_fu_arch_n510) );
  AOI22X2 fu_ALU_fu_arch_U194 ( .A0(n2100), .A1(n1882), .B0(
        fu_ALU_fu_arch_n333), .B1(fu_ALU_fu_arch_n345), .Y(fu_ALU_fu_arch_n419) );
  AOI22X2 fu_ALU_fu_arch_U281 ( .A0(fu_ALU_fu_arch_n333), .A1(n1795), .B0(
        n2101), .B1(n1838), .Y(fu_ALU_fu_arch_n521) );
  AOI22X2 U443 ( .A0(ic_socket_gcu_o1_data0_wire[11]), .A1(n2115), .B0(n2116), 
        .B1(inst_fetch_increased_pc_11_), .Y(n299) );
  AOI22X2 fu_ALU_fu_arch_U211 ( .A0(n2100), .A1(n1795), .B0(
        fu_ALU_fu_arch_n333), .B1(fu_ALU_fu_arch_n366), .Y(fu_ALU_fu_arch_n443) );
  INVX2 U799 ( .A(n448), .Y(n447) );
  AOI222X2 fu_ALU_fu_arch_U216 ( .A0(fu_ALU_o1reg[24]), .A1(
        fu_ALU_fu_arch_n450), .B0(n2101), .B1(n1840), .C0(fu_ALU_fu_arch_n395), 
        .C1(n1838), .Y(fu_ALU_fu_arch_n449) );
  AOI22X2 fu_ALU_fu_arch_U413 ( .A0(n2103), .A1(n1836), .B0(n1892), .B1(n1835), 
        .Y(fu_ALU_fu_arch_n642) );
  AOI22X2 fu_ALU_fu_arch_U199 ( .A0(n2101), .A1(n1796), .B0(
        fu_ALU_fu_arch_n395), .B1(n1845), .Y(fu_ALU_fu_arch_n427) );
  AOI22X2 fu_ALU_fu_arch_U432 ( .A0(n2103), .A1(fu_ALU_fu_arch_n435), .B0(
        n2156), .B1(fu_ALU_fu_arch_n153), .Y(fu_ALU_fu_arch_n657) );
  NAND2X2 fu_ALU_fu_arch_U223 ( .A(fu_ALU_fu_arch_n147), .B(
        fu_ALU_fu_arch_n437), .Y(fu_ALU_fu_arch_n142) );
  AOI22X2 U791 ( .A0(ic_socket_lsu_o1_data0_wire[6]), .A1(n2212), .B0(n1280), 
        .B1(fu_LSU_data_in[22]), .Y(n444) );
  AOI22X2 fu_ALU_fu_arch_U527 ( .A0(n1854), .A1(n1834), .B0(
        fu_ALU_fu_arch_n178), .B1(fu_ALU_fu_arch_n399), .Y(fu_ALU_fu_arch_n693) );
  AOI22X2 U784 ( .A0(ic_socket_lsu_o1_data0_wire[4]), .A1(n2212), .B0(n1280), 
        .B1(fu_LSU_data_in[20]), .Y(n438) );
  AOI22X2 U787 ( .A0(ic_socket_lsu_o1_data0_wire[5]), .A1(n2212), .B0(n1280), 
        .B1(fu_LSU_data_in[21]), .Y(n441) );
  OAI21X4 fu_ALU_fu_arch_U248 ( .A0(n1807), .A1(fu_ALU_fu_arch_n468), .B0(
        fu_ALU_fu_arch_n488), .Y(fu_ALU_fu_arch_n191) );
  AOI22X2 U775 ( .A0(ic_socket_lsu_o1_data0_wire[1]), .A1(n2212), .B0(n1280), 
        .B1(fu_LSU_data_in[17]), .Y(n429) );
  AOI22X2 U781 ( .A0(ic_socket_lsu_o1_data0_wire[3]), .A1(n2212), .B0(n1280), 
        .B1(fu_LSU_data_in[19]), .Y(n435) );
  NAND2X2 fu_ALU_fu_arch_U405 ( .A(fu_ALU_fu_arch_n637), .B(
        fu_ALU_fu_arch_n638), .Y(fu_ALU_fu_arch_n277) );
  AOI211X4 fu_ALU_fu_arch_U83 ( .A0(n2174), .A1(fu_ALU_fu_arch_n169), .B0(
        fu_ALU_fu_arch_n232), .C0(fu_ALU_fu_arch_n233), .Y(fu_ALU_fu_arch_n231) );
  AOI22X2 fu_ALU_fu_arch_U228 ( .A0(fu_ALU_fu_arch_n240), .A1(
        fu_ALU_fu_arch_n179), .B0(fu_ALU_fu_arch_n333), .B1(n1793), .Y(
        fu_ALU_fu_arch_n465) );
  AOI32X2 fu_ALU_fu_arch_U119 ( .A0(n1850), .A1(fu_ALU_fu_arch_n304), .A2(
        n2172), .B0(fu_ALU_fu_arch_n305), .B1(n1850), .Y(fu_ALU_fu_arch_n293)
         );
  AOI22X2 fu_ALU_fu_arch_U565 ( .A0(fu_ALU_fu_arch_n111), .A1(
        fu_ALU_fu_arch_n405), .B0(fu_ALU_fu_arch_n178), .B1(
        fu_ALU_fu_arch_n416), .Y(fu_ALU_fu_arch_n717) );
  AOI22X2 U778 ( .A0(ic_socket_lsu_o1_data0_wire[2]), .A1(n2212), .B0(n1280), 
        .B1(fu_LSU_data_in[18]), .Y(n432) );
  OAI211X2 fu_ALU_fu_arch_U170 ( .A0(fu_ALU_fu_arch_n387), .A1(
        fu_ALU_fu_arch_n388), .B0(fu_ALU_fu_arch_n389), .C0(
        fu_ALU_fu_arch_n390), .Y(fu_ALU_fu_arch_n386) );
  AOI22X2 fu_ALU_fu_arch_U37 ( .A0(n2191), .A1(fu_ALU_fu_arch_N620), .B0(n2193), .B1(fu_ALU_fu_arch_N41), .Y(fu_ALU_fu_arch_n151) );
  AOI222X2 U821 ( .A0(ic_socket_lsu_o1_data0_wire[15]), .A1(n2212), .B0(n457), 
        .B1(n474), .C0(n2118), .C1(fu_LSU_data_in[15]), .Y(n473) );
  AOI22X2 fu_ALU_fu_arch_U154 ( .A0(n2172), .A1(fu_ALU_fu_arch_n364), .B0(
        fu_ALU_fu_arch_n365), .B1(fu_ALU_fu_arch_n220), .Y(fu_ALU_fu_arch_n363) );
  NAND2X2 fu_ALU_fu_arch_U233 ( .A(fu_ALU_fu_arch_n472), .B(n2102), .Y(
        fu_ALU_fu_arch_n471) );
  AOI22X2 U772 ( .A0(ic_socket_lsu_o1_data0_wire[0]), .A1(n2212), .B0(n1280), 
        .B1(fu_LSU_data_in[16]), .Y(n422) );
  AOI22X2 U414 ( .A0(ic_socket_gcu_o1_data0_wire[12]), .A1(n2115), .B0(n2116), 
        .B1(inst_fetch_increased_pc_12_), .Y(n288) );
  NAND2X2 fu_ALU_fu_arch_U207 ( .A(fu_ALU_fu_arch_n436), .B(
        fu_ALU_fu_arch_n437), .Y(fu_ALU_fu_arch_n112) );
  OAI211X2 fu_ALU_fu_arch_U198 ( .A0(fu_ALU_fu_arch_n425), .A1(n2134), .B0(
        fu_ALU_fu_arch_n427), .C0(n2102), .Y(fu_ALU_fu_arch_n424) );
  AOI22X2 U402 ( .A0(busy), .A1(inst_fetch_pc_reg_12_), .B0(n2114), .B1(
        inst_fetch_increased_pc_12_), .Y(n287) );
  NAND2X2 fu_ALU_fu_arch_U285 ( .A(fu_ALU_fu_arch_n527), .B(n2102), .Y(
        fu_ALU_fu_arch_n526) );
  NAND2X2 fu_ALU_fu_arch_U215 ( .A(fu_ALU_fu_arch_n449), .B(n2102), .Y(
        fu_ALU_fu_arch_n448) );
  AOI22X2 U373 ( .A0(busy), .A1(inst_fetch_pc_reg_13_), .B0(n2114), .B1(
        inst_fetch_increased_pc_13_), .Y(n274) );
  NOR2X2 U752 ( .A(n2185), .B(n2249), .Y(n219) );
  AOI22X2 fu_ALU_fu_arch_U245 ( .A0(fu_ALU_fu_arch_n240), .A1(
        fu_ALU_fu_arch_n191), .B0(fu_ALU_fu_arch_n333), .B1(n1794), .Y(
        fu_ALU_fu_arch_n485) );
  NAND2X2 fu_ALU_fu_arch_U11 ( .A(fu_ALU_fu_arch_n111), .B(fu_ALU_fu_arch_n112), .Y(fu_ALU_fu_arch_n110) );
  AOI22X2 fu_ALU_fu_arch_U141 ( .A0(n2172), .A1(fu_ALU_fu_arch_n343), .B0(
        fu_ALU_fu_arch_n344), .B1(fu_ALU_fu_arch_n220), .Y(fu_ALU_fu_arch_n342) );
  AOI22X2 fu_ALU_fu_arch_U103 ( .A0(n2172), .A1(fu_ALU_fu_arch_n277), .B0(
        fu_ALU_fu_arch_n278), .B1(fu_ALU_fu_arch_n279), .Y(fu_ALU_fu_arch_n276) );
  AOI22X2 U385 ( .A0(ic_socket_gcu_o1_data0_wire[13]), .A1(n2115), .B0(n2116), 
        .B1(inst_fetch_increased_pc_13_), .Y(n277) );
  AOI22X2 U363 ( .A0(ic_socket_gcu_o1_data0_wire[14]), .A1(n2115), .B0(
        inst_fetch_increased_pc_14_), .B1(n2116), .Y(n265) );
  AOI22X2 fu_ALU_fu_arch_U549 ( .A0(n2191), .A1(fu_ALU_fu_arch_N622), .B0(
        n2194), .B1(fu_ALU_fu_arch_N43), .Y(fu_ALU_fu_arch_n722) );
  AOI22X2 U910 ( .A0(busy), .A1(inst_fetch_pc_reg_14_), .B0(
        inst_fetch_increased_pc_14_), .B1(n2114), .Y(n506) );
  NAND2X2 U314 ( .A(n2120), .B(fu_LSU_o1shadow_reg_16_), .Y(n237) );
  AOI22X2 U815 ( .A0(fu_LSU_data_in[14]), .A1(n1863), .B0(
        ic_socket_lsu_o1_data0_wire[14]), .B1(n2212), .Y(n469) );
  AOI22X2 U248 ( .A0(fu_LSU_o1shadow_reg_19_), .A1(n2120), .B0(
        fu_LSU_data_out[19]), .B1(n2248), .Y(n192) );
  AOI22X2 U206 ( .A0(fu_LSU_o1shadow_reg_21_), .A1(n2120), .B0(
        fu_LSU_data_out[21]), .B1(n2248), .Y(n168) );
  AOI22X2 U813 ( .A0(fu_LSU_data_in[13]), .A1(n1863), .B0(
        ic_socket_lsu_o1_data0_wire[13]), .B1(n2212), .Y(n468) );
  AOI22X2 U227 ( .A0(fu_LSU_o1shadow_reg_20_), .A1(n2120), .B0(
        fu_LSU_data_out[20]), .B1(n2248), .Y(n180) );
  AOI22X2 U185 ( .A0(fu_LSU_o1shadow_reg_22_), .A1(n2120), .B0(
        fu_LSU_data_out[22]), .B1(n2248), .Y(n156) );
  AOI22X2 U811 ( .A0(fu_LSU_data_in[12]), .A1(n1863), .B0(
        ic_socket_lsu_o1_data0_wire[12]), .B1(n2212), .Y(n467) );
  AOI22X2 U95 ( .A0(fu_LSU_o1shadow_reg_26_), .A1(n2120), .B0(
        fu_LSU_data_out[26]), .B1(n2249), .Y(n100) );
  OAI211X2 fu_ALU_fu_arch_U548 ( .A0(fu_ALU_fu_arch_n408), .A1(
        fu_ALU_fu_arch_n108), .B0(fu_ALU_fu_arch_n721), .C0(
        fu_ALU_fu_arch_n722), .Y(fu_ALU_fu_arch_n720) );
  AOI22X2 U269 ( .A0(fu_LSU_o1shadow_reg_18_), .A1(n2120), .B0(
        fu_LSU_data_out[18]), .B1(n2248), .Y(n204) );
  AOI22X2 U73 ( .A0(fu_LSU_o1shadow_reg_27_), .A1(n2120), .B0(
        fu_LSU_data_out[27]), .B1(n2249), .Y(n88) );
  AOI22X2 U10 ( .A0(fu_LSU_o1shadow_reg_30_), .A1(n2120), .B0(
        fu_LSU_data_out[30]), .B1(n2249), .Y(n36) );
  NAND2X2 U751 ( .A(fu_LSU_o1shadow_reg_0_), .B(n2121), .Y(n235) );
  AOI22X2 U805 ( .A0(fu_LSU_data_in[9]), .A1(n1863), .B0(
        ic_socket_lsu_o1_data0_wire[9]), .B1(n2212), .Y(n464) );
  AOI22X2 U807 ( .A0(fu_LSU_data_in[10]), .A1(n1863), .B0(
        ic_socket_lsu_o1_data0_wire[10]), .B1(n2212), .Y(n465) );
  AOI22X2 U803 ( .A0(fu_LSU_data_in[8]), .A1(n1863), .B0(
        ic_socket_lsu_o1_data0_wire[8]), .B1(n2212), .Y(n461) );
  AOI22X2 U290 ( .A0(fu_LSU_o1shadow_reg_17_), .A1(n2120), .B0(
        fu_LSU_data_out[17]), .B1(n2248), .Y(n218) );
  AOI22X2 U31 ( .A0(fu_LSU_o1shadow_reg_29_), .A1(n2120), .B0(
        fu_LSU_data_out[29]), .B1(n2249), .Y(n63) );
  AOI22X2 U52 ( .A0(fu_LSU_o1shadow_reg_28_), .A1(n2120), .B0(
        fu_LSU_data_out[28]), .B1(n2248), .Y(n76) );
  AOI22X2 U5 ( .A0(fu_LSU_o1shadow_reg_31_), .A1(n2120), .B0(
        fu_LSU_data_out[31]), .B1(n2249), .Y(n26) );
  AOI22X2 U139 ( .A0(fu_LSU_o1shadow_reg_24_), .A1(n2120), .B0(
        fu_LSU_data_out[24]), .B1(n2248), .Y(n126) );
  AOI22X2 fu_ALU_fu_arch_U504 ( .A0(n2192), .A1(fu_ALU_fu_arch_N623), .B0(
        n2194), .B1(fu_ALU_fu_arch_N44), .Y(fu_ALU_fu_arch_n699) );
  AOI22X2 U762 ( .A0(fu_LSU_o1shadow_reg_1_), .A1(n2120), .B0(
        fu_LSU_data_out[1]), .B1(n2248), .Y(n414) );
  AOI22X2 U117 ( .A0(fu_LSU_o1shadow_reg_25_), .A1(n2120), .B0(
        fu_LSU_data_out[25]), .B1(n2249), .Y(n116) );
  AOI22X2 U164 ( .A0(fu_LSU_o1shadow_reg_23_), .A1(n2120), .B0(
        fu_LSU_data_out[23]), .B1(n2248), .Y(n143) );
  AOI22X2 fu_ALU_fu_arch_U99 ( .A0(n1850), .A1(fu_ALU_fu_arch_n267), .B0(
        fu_ALU_o1reg[31]), .B1(fu_ALU_fu_arch_n268), .Y(fu_ALU_fu_arch_n265)
         );
  AOI22X2 U809 ( .A0(fu_LSU_data_in[11]), .A1(n1863), .B0(
        ic_socket_lsu_o1_data0_wire[11]), .B1(n2212), .Y(n466) );
  OAI211X2 fu_ALU_fu_arch_U29 ( .A0(fu_ALU_fu_arch_n139), .A1(
        fu_ALU_fu_arch_n108), .B0(fu_ALU_fu_arch_n140), .C0(
        fu_ALU_fu_arch_n141), .Y(ic_socket_ALU_o1_data0_wire[8]) );
  AOI22X2 U774 ( .A0(fu_LSU_data_in[9]), .A1(n1858), .B0(fu_LSU_data_in[1]), 
        .B1(n1287), .Y(n430) );
  OAI211X2 U806 ( .A0(n431), .A1(n460), .B0(n465), .C0(n462), .Y(n1043) );
  OAI211X2 U802 ( .A0(n421), .A1(n460), .B0(n461), .C0(n462), .Y(n1041) );
  AOI22X2 U777 ( .A0(fu_LSU_data_in[10]), .A1(n1858), .B0(fu_LSU_data_in[2]), 
        .B1(n1287), .Y(n433) );
  OAI211X2 U804 ( .A0(n428), .A1(n460), .B0(n464), .C0(n462), .Y(n1042) );
  AOI22X2 U789 ( .A0(fu_LSU_data_in[14]), .A1(n1858), .B0(fu_LSU_data_in[6]), 
        .B1(n1287), .Y(n445) );
  AOI22X2 U771 ( .A0(fu_LSU_data_in[8]), .A1(n1858), .B0(fu_LSU_data_in[0]), 
        .B1(n1287), .Y(n423) );
  NAND2BX2 U820 ( .AN(n2119), .B(n473), .Y(n1048) );
  AOI22X2 fu_ALU_fu_arch_U486 ( .A0(n2192), .A1(fu_ALU_fu_arch_N624), .B0(
        n2194), .B1(fu_ALU_fu_arch_N45), .Y(fu_ALU_fu_arch_n685) );
  AOI22X2 U786 ( .A0(fu_LSU_data_in[13]), .A1(n1858), .B0(fu_LSU_data_in[5]), 
        .B1(n1287), .Y(n442) );
  AOI22X2 U780 ( .A0(fu_LSU_data_in[11]), .A1(n1858), .B0(fu_LSU_data_in[3]), 
        .B1(n1287), .Y(n436) );
  AOI22X2 U783 ( .A0(fu_LSU_data_in[12]), .A1(n1858), .B0(fu_LSU_data_in[4]), 
        .B1(n1287), .Y(n439) );
  OAI211X2 U810 ( .A0(n437), .A1(n460), .B0(n467), .C0(n462), .Y(n1045) );
  OAI211X2 U808 ( .A0(n434), .A1(n460), .B0(n466), .C0(n462), .Y(n1044) );
  AOI22X2 U795 ( .A0(fu_LSU_data_in[23]), .A1(n1280), .B0(fu_LSU_data_in[7]), 
        .B1(n1287), .Y(n450) );
  OAI211X2 U812 ( .A0(n440), .A1(n460), .B0(n468), .C0(n462), .Y(n1046) );
  OAI211X2 fu_ALU_fu_arch_U503 ( .A0(fu_ALU_fu_arch_n387), .A1(
        fu_ALU_fu_arch_n108), .B0(fu_ALU_fu_arch_n698), .C0(
        fu_ALU_fu_arch_n699), .Y(fu_ALU_fu_arch_n697) );
  OAI211X2 U814 ( .A0(n443), .A1(n460), .B0(n469), .C0(n462), .Y(n1047) );
  OAI211X2 fu_ALU_fu_arch_U10 ( .A0(fu_ALU_fu_arch_n107), .A1(
        fu_ALU_fu_arch_n108), .B0(fu_ALU_fu_arch_n109), .C0(
        fu_ALU_fu_arch_n110), .Y(ic_socket_ALU_o1_data0_wire[9]) );
  OAI211X2 U788 ( .A0(n420), .A1(n443), .B0(n444), .C0(n445), .Y(n1039) );
  OAI211X2 U793 ( .A0(n1806), .A1(n447), .B0(n450), .C0(n451), .Y(n1040) );
  OAI211X2 fu_ALU_fu_arch_U62 ( .A0(fu_ALU_fu_arch_n131), .A1(
        fu_ALU_fu_arch_n136), .B0(fu_ALU_fu_arch_n196), .C0(
        fu_ALU_fu_arch_n197), .Y(ic_socket_ALU_o1_data0_wire[5]) );
  AOI22X2 fu_ALU_fu_arch_U439 ( .A0(n2192), .A1(fu_ALU_fu_arch_N625), .B0(
        n2194), .B1(fu_ALU_fu_arch_N46), .Y(fu_ALU_fu_arch_n662) );
  OAI211X2 U773 ( .A0(n420), .A1(n428), .B0(n429), .C0(n430), .Y(n1034) );
  OAI211X2 U770 ( .A0(n420), .A1(n421), .B0(n422), .C0(n423), .Y(n1033) );
  OAI211X2 U785 ( .A0(n420), .A1(n440), .B0(n441), .C0(n442), .Y(n1038) );
  OAI211X2 U782 ( .A0(n420), .A1(n437), .B0(n438), .C0(n439), .Y(n1037) );
  OAI211X2 U779 ( .A0(n420), .A1(n434), .B0(n435), .C0(n436), .Y(n1036) );
  OAI211X2 U776 ( .A0(n420), .A1(n431), .B0(n432), .C0(n433), .Y(n1035) );
  AOI22X2 U566 ( .A0(fu_ALU_o1reg[6]), .A1(n2252), .B0(n2251), .B1(n1818), .Y(
        n354) );
  AOI22X2 U620 ( .A0(fu_ALU_fu_arch_sub_200_B_4_), .A1(n2253), .B0(n2250), 
        .B1(n1825), .Y(n374) );
  AOI22X2 U539 ( .A0(n2166), .A1(n2253), .B0(n2251), .B1(n1814), .Y(n343) );
  AOI22X2 fu_ALU_fu_arch_U424 ( .A0(n2192), .A1(fu_ALU_fu_arch_N626), .B0(
        n2193), .B1(fu_ALU_fu_arch_N47), .Y(fu_ALU_fu_arch_n649) );
  OAI211X2 fu_ALU_fu_arch_U437 ( .A0(fu_ALU_fu_arch_n343), .A1(
        fu_ALU_fu_arch_n108), .B0(fu_ALU_fu_arch_n662), .C0(
        fu_ALU_fu_arch_n663), .Y(fu_ALU_fu_arch_n661) );
  INVX2 U397 ( .A(n179), .Y(n78) );
  AOI2BB2X2 U581 ( .B0(n2227), .B1(n355), .A0N(rf_RF_reg_3__6_), .A1N(n2229), 
        .Y(n930) );
  AOI2BB2X2 U890 ( .B0(n2235), .B1(n2117), .A0N(rf_RF_reg_1__1_), .A1N(n2238), 
        .Y(n1069) );
  AOI2BB2X2 U892 ( .B0(n2227), .B1(n2117), .A0N(rf_RF_reg_3__1_), .A1N(n2230), 
        .Y(n1071) );
  AOI22X2 U630 ( .A0(n1285), .A1(n375), .B0(n373), .B1(n2244), .Y(n956) );
  AOI2BB2X2 U893 ( .B0(n2223), .B1(n2117), .A0N(rf_RF_reg_4__1_), .A1N(n2226), 
        .Y(n1072) );
  AOI2BB2X2 U891 ( .B0(n2231), .B1(n2117), .A0N(rf_RF_reg_2__1_), .A1N(n2234), 
        .Y(n1070) );
  AOI2BB2X2 U580 ( .B0(n2231), .B1(n355), .A0N(rf_RF_reg_2__6_), .A1N(n2233), 
        .Y(n929) );
  AOI2BB2X2 U578 ( .B0(n2239), .B1(n355), .A0N(rf_RF_reg_0__6_), .A1N(n2241), 
        .Y(n927) );
  AOI2BB2X2 U553 ( .B0(n2231), .B1(n345), .A0N(rf_RF_reg_2__7_), .A1N(n2233), 
        .Y(n914) );
  AOI2BB2X2 U551 ( .B0(n2239), .B1(n345), .A0N(rf_RF_reg_0__7_), .A1N(n2241), 
        .Y(n912) );
  OAI211X2 fu_ALU_fu_arch_U477 ( .A0(fu_ALU_fu_arch_n364), .A1(
        fu_ALU_fu_arch_n108), .B0(fu_ALU_fu_arch_n676), .C0(
        fu_ALU_fu_arch_n677), .Y(ic_socket_ALU_o1_data0_wire[12]) );
  AOI2BB2X2 U582 ( .B0(n2223), .B1(n355), .A0N(rf_RF_reg_4__6_), .A1N(n2225), 
        .Y(n931) );
  AOI2BB2X2 U579 ( .B0(n2235), .B1(n355), .A0N(rf_RF_reg_1__6_), .A1N(n2237), 
        .Y(n928) );
  AOI2BB2X2 U889 ( .B0(n2239), .B1(n2117), .A0N(rf_RF_reg_0__1_), .A1N(n2242), 
        .Y(n1068) );
  AOI2BB2X2 U555 ( .B0(n2223), .B1(n345), .A0N(rf_RF_reg_4__7_), .A1N(n2225), 
        .Y(n916) );
  AOI2BB2X2 U554 ( .B0(n2227), .B1(n345), .A0N(rf_RF_reg_3__7_), .A1N(n2229), 
        .Y(n915) );
  AOI2BB2X2 U552 ( .B0(n2235), .B1(n345), .A0N(rf_RF_reg_1__7_), .A1N(n2237), 
        .Y(n913) );
  AOI2BB2X2 U632 ( .B0(n2239), .B1(n375), .A0N(rf_RF_reg_0__4_), .A1N(n2242), 
        .Y(n957) );
  AOI2BB2X2 U634 ( .B0(n2231), .B1(n375), .A0N(rf_RF_reg_2__4_), .A1N(n2234), 
        .Y(n959) );
  INVX2 U360 ( .A(n155), .Y(n38) );
  AOI2BB2X2 U628 ( .B0(n2245), .B1(n375), .A0N(fu_LSU_o1shadow_reg_4_), .A1N(
        n2246), .Y(n954) );
  AOI2BB2X2 U636 ( .B0(n2223), .B1(n375), .A0N(rf_RF_reg_4__4_), .A1N(n2226), 
        .Y(n961) );
  AOI22X2 U768 ( .A0(n2245), .A1(n2117), .B0(n115), .B1(n419), .Y(n1032) );
  AOI2BB2X2 U635 ( .B0(n2227), .B1(n375), .A0N(rf_RF_reg_3__4_), .A1N(n2230), 
        .Y(n960) );
  AOI2BB2X2 U633 ( .B0(n2235), .B1(n375), .A0N(rf_RF_reg_1__4_), .A1N(n2238), 
        .Y(n958) );
  NAND3X2 fu_ALU_fu_arch_U419 ( .A(fu_ALU_fu_arch_n649), .B(
        fu_ALU_fu_arch_n650), .C(fu_ALU_fu_arch_n651), .Y(fu_ALU_fu_arch_n643)
         );
  INVX2 U338 ( .A(n141), .Y(n30) );
  AOI22X2 U703 ( .A0(n2177), .A1(n2253), .B0(n2250), .B1(n2110), .Y(n404) );
  AOI22X2 U549 ( .A0(n1285), .A1(n345), .B0(n342), .B1(n2244), .Y(n911) );
  AOI22X2 U885 ( .A0(n500), .A1(n2117), .B0(n499), .B1(n501), .Y(n1066) );
  AOI2BB2X2 U574 ( .B0(n2245), .B1(n355), .A0N(fu_LSU_o1shadow_reg_6_), .A1N(
        n2246), .Y(n924) );
  AOI22X2 U887 ( .A0(n1761), .A1(n2117), .B0(n403), .B1(n2243), .Y(n1067) );
  AOI22X2 U647 ( .A0(n2173), .A1(n2253), .B0(n2251), .B1(n1808), .Y(n384) );
  AOI22X2 U674 ( .A0(fu_ALU_fu_arch_sub_200_B_2_), .A1(n2253), .B0(n2250), 
        .B1(n1810), .Y(n394) );
  AOI22X2 U576 ( .A0(n1285), .A1(n355), .B0(n353), .B1(n2244), .Y(n926) );
  AOI2BB2X2 U547 ( .B0(n2245), .B1(n345), .A0N(fu_LSU_o1shadow_reg_7_), .A1N(
        n2246), .Y(n909) );
  AOI22X2 U657 ( .A0(n1761), .A1(n385), .B0(n383), .B1(n2243), .Y(n971) );
  INVX2 U426 ( .A(n191), .Y(n90) );
  AOI2BB2X2 U691 ( .B0(n2227), .B1(n395), .A0N(rf_RF_reg_3__2_), .A1N(n2230), 
        .Y(n990) );
  AOI2BB2X2 U660 ( .B0(n2235), .B1(n385), .A0N(rf_RF_reg_1__3_), .A1N(n2238), 
        .Y(n973) );
  AOI2BB2X2 U659 ( .B0(n2239), .B1(n385), .A0N(rf_RF_reg_0__3_), .A1N(n2242), 
        .Y(n972) );
  AOI2BB2X2 U662 ( .B0(n2227), .B1(n385), .A0N(rf_RF_reg_3__3_), .A1N(n2230), 
        .Y(n975) );
  AOI2BB2X2 U689 ( .B0(n2235), .B1(n395), .A0N(rf_RF_reg_1__2_), .A1N(n2238), 
        .Y(n988) );
  AOI22X2 U686 ( .A0(n1761), .A1(n395), .B0(n393), .B1(n2244), .Y(n986) );
  AOI2BB2X2 U661 ( .B0(n2231), .B1(n385), .A0N(rf_RF_reg_2__3_), .A1N(n2234), 
        .Y(n974) );
  AOI2BB2X2 U692 ( .B0(n2223), .B1(n395), .A0N(rf_RF_reg_4__2_), .A1N(n2226), 
        .Y(n991) );
  AOI2BB2X2 U688 ( .B0(n2239), .B1(n395), .A0N(rf_RF_reg_0__2_), .A1N(n2242), 
        .Y(n987) );
  AOI2BB2X2 U690 ( .B0(n2231), .B1(n395), .A0N(rf_RF_reg_2__2_), .A1N(n2234), 
        .Y(n989) );
  AOI2BB2X2 U528 ( .B0(n2223), .B1(n2122), .A0N(rf_RF_reg_4__8_), .A1N(n2226), 
        .Y(n901) );
  INVX2 U138 ( .A(n25), .Y(n128) );
  AOI2BB2X2 U663 ( .B0(n2223), .B1(n385), .A0N(rf_RF_reg_4__3_), .A1N(n2226), 
        .Y(n976) );
  AOI2BB2X2 U525 ( .B0(n2235), .B1(n2122), .A0N(rf_RF_reg_1__8_), .A1N(n2238), 
        .Y(n898) );
  AOI2BB2X2 U526 ( .B0(n2231), .B1(n2122), .A0N(rf_RF_reg_2__8_), .A1N(n2234), 
        .Y(n899) );
  AOI2BB2X2 U524 ( .B0(n2239), .B1(n2122), .A0N(rf_RF_reg_0__8_), .A1N(n2242), 
        .Y(n897) );
  AOI22X2 U522 ( .A0(n1285), .A1(n2122), .B0(n329), .B1(n2244), .Y(n896) );
  INVX2 U455 ( .A(n203), .Y(n102) );
  AOI2BB2X2 U655 ( .B0(n2245), .B1(n385), .A0N(fu_LSU_o1shadow_reg_3_), .A1N(
        n2245), .Y(n969) );
  AOI22X2 U481 ( .A0(fu_ALU_fu_arch_sub_200_B_9_), .A1(n2253), .B0(n2251), 
        .B1(n1812), .Y(n317) );
  AOI2BB2X2 U684 ( .B0(n2245), .B1(n395), .A0N(fu_LSU_o1shadow_reg_2_), .A1N(
        n2245), .Y(n984) );
  OAI2B11X2 fu_ALU_fu_arch_U431 ( .A1N(fu_ALU_fu_arch_n636), .A0(
        fu_ALU_fu_arch_n337), .B0(fu_ALU_fu_arch_n656), .C0(
        fu_ALU_fu_arch_n657), .Y(ic_socket_ALU_o1_data0_wire[13]) );
  AOI2BB2X2 U520 ( .B0(n2245), .B1(n2122), .A0N(fu_LSU_o1shadow_reg_8_), .A1N(
        n2246), .Y(n894) );
  AOI2BB2X2 U527 ( .B0(n2227), .B1(n2122), .A0N(rf_RF_reg_3__8_), .A1N(n2230), 
        .Y(n900) );
  AOI22X2 U452 ( .A0(n2161), .A1(n2252), .B0(n2251), .B1(n1816), .Y(n306) );
  AOI22X2 U593 ( .A0(fu_ALU_o1reg[5]), .A1(n2253), .B0(n2250), .B1(n1821), .Y(
        n364) );
  AOI22X2 U493 ( .A0(n1285), .A1(n321), .B0(n316), .B1(n2244), .Y(n881) );
  AOI2BB2X2 U491 ( .B0(n2245), .B1(n321), .A0N(fu_LSU_o1shadow_reg_9_), .A1N(
        n2246), .Y(n879) );
  NAND3X2 fu_ALU_fu_arch_U412 ( .A(fu_ALU_fu_arch_n640), .B(
        fu_ALU_fu_arch_n641), .C(fu_ALU_fu_arch_n642), .Y(
        ic_socket_ALU_o1_data0_wire[14]) );
  AOI2BB2X2 U497 ( .B0(n2231), .B1(n321), .A0N(rf_RF_reg_2__9_), .A1N(n2233), 
        .Y(n884) );
  AOI2BB2X2 U496 ( .B0(n2235), .B1(n321), .A0N(rf_RF_reg_1__9_), .A1N(n2237), 
        .Y(n883) );
  AOI22X2 fu_ALU_fu_arch_U363 ( .A0(n2192), .A1(fu_ALU_fu_arch_N629), .B0(
        n2193), .B1(fu_ALU_fu_arch_N50), .Y(fu_ALU_fu_arch_n603) );
  AOI2BB2X2 U495 ( .B0(n2239), .B1(n321), .A0N(rf_RF_reg_0__9_), .A1N(n2241), 
        .Y(n882) );
  AOI2BB2X2 U499 ( .B0(n2223), .B1(n321), .A0N(rf_RF_reg_4__9_), .A1N(n2225), 
        .Y(n886) );
  NAND2X2 U1142 ( .A(n601), .B(n2111), .Y(n557) );
  AOI2BB2X2 U498 ( .B0(n2227), .B1(n321), .A0N(rf_RF_reg_3__9_), .A1N(n2229), 
        .Y(n885) );
  AOI2BB2X2 U470 ( .B0(n2223), .B1(n308), .A0N(rf_RF_reg_4__10_), .A1N(n2225), 
        .Y(n871) );
  AOI2BB2X2 U467 ( .B0(n2235), .B1(n308), .A0N(rf_RF_reg_1__10_), .A1N(n2237), 
        .Y(n868) );
  AOI2BB2X2 U466 ( .B0(n2239), .B1(n308), .A0N(rf_RF_reg_0__10_), .A1N(n2241), 
        .Y(n867) );
  AOI2BB2X2 U469 ( .B0(n2227), .B1(n308), .A0N(rf_RF_reg_3__10_), .A1N(n2229), 
        .Y(n870) );
  OAI211X2 fu_ALU_fu_arch_U362 ( .A0(fu_ALU_fu_arch_n510), .A1(
        fu_ALU_fu_arch_n235), .B0(fu_ALU_fu_arch_n602), .C0(
        fu_ALU_fu_arch_n603), .Y(fu_ALU_fu_arch_n599) );
  AOI2BB2X2 U605 ( .B0(n2239), .B1(n365), .A0N(rf_RF_reg_0__5_), .A1N(n2242), 
        .Y(n942) );
  AOI22X2 fu_ALU_fu_arch_U344 ( .A0(n2192), .A1(fu_ALU_fu_arch_N630), .B0(
        n2193), .B1(fu_ALU_fu_arch_N51), .Y(fu_ALU_fu_arch_n587) );
  AOI2BB2X2 U607 ( .B0(n2231), .B1(n365), .A0N(rf_RF_reg_2__5_), .A1N(n2234), 
        .Y(n944) );
  NAND3X2 fu_ALU_fu_arch_U394 ( .A(fu_ALU_fu_arch_n624), .B(
        fu_ALU_fu_arch_n625), .C(fu_ALU_fu_arch_n626), .Y(
        ic_socket_ALU_o1_data0_wire[15]) );
  AOI2BB2X2 U468 ( .B0(n2231), .B1(n308), .A0N(rf_RF_reg_2__10_), .A1N(n2233), 
        .Y(n869) );
  NAND3X2 U1145 ( .A(inst_decoder_instructionword_wire[41]), .B(n597), .C(n603), .Y(n593) );
  AOI22X2 U512 ( .A0(n332), .A1(n129), .B0(fu_LSU_data_out[8]), .B1(n2248), 
        .Y(n331) );
  INVX2 U368 ( .A(n167), .Y(n65) );
  AOI2BB2X2 U462 ( .B0(n2245), .B1(n308), .A0N(fu_LSU_o1shadow_reg_10_), .A1N(
        n2246), .Y(n864) );
  AOI2BB2X2 U601 ( .B0(n2245), .B1(n365), .A0N(fu_LSU_o1shadow_reg_5_), .A1N(
        n2246), .Y(n939) );
  AOI2BB2X2 U609 ( .B0(n2223), .B1(n365), .A0N(rf_RF_reg_4__5_), .A1N(n2226), 
        .Y(n946) );
  AOI22X2 U464 ( .A0(n1285), .A1(n308), .B0(n305), .B1(n2244), .Y(n866) );
  AOI2BB2X2 U606 ( .B0(n2235), .B1(n365), .A0N(rf_RF_reg_1__5_), .A1N(n2238), 
        .Y(n943) );
  AOI2BB2X2 U608 ( .B0(n2227), .B1(n365), .A0N(rf_RF_reg_3__5_), .A1N(n2230), 
        .Y(n945) );
  AOI22X2 fu_ALU_fu_arch_U290 ( .A0(n2193), .A1(fu_ALU_fu_arch_N53), .B0(n2145), .B1(fu_ALU_fu_arch_n532), .Y(fu_ALU_fu_arch_n531) );
  NAND2X2 U1138 ( .A(n220), .B(n601), .Y(n600) );
  AOI22X2 U351 ( .A0(n2257), .A1(ic_socket_ALU_o1_data0_wire[15]), .B0(n2222), 
        .B1(rf_RF_reg_4__15_), .Y(n256) );
  AOI22X2 fu_ALU_fu_arch_U325 ( .A0(n2192), .A1(fu_ALU_fu_arch_N631), .B0(
        n2193), .B1(fu_ALU_fu_arch_N52), .Y(fu_ALU_fu_arch_n570) );
  NAND2X2 U514 ( .A(n1270), .B(n2110), .Y(n320) );
  OAI211X2 fu_ALU_fu_arch_U343 ( .A0(fu_ALU_fu_arch_n483), .A1(
        fu_ALU_fu_arch_n235), .B0(fu_ALU_fu_arch_n586), .C0(
        fu_ALU_fu_arch_n587), .Y(fu_ALU_fu_arch_n584) );
  AOI22X2 U423 ( .A0(fu_ALU_fu_arch_sub_200_B_11_), .A1(n2253), .B0(n2251), 
        .B1(rf_RF_t1data_wire[11]), .Y(n295) );
  AOI2BB2X2 U433 ( .B0(n2245), .B1(n297), .A0N(fu_LSU_o1shadow_reg_11_), .A1N(
        n2246), .Y(n849) );
  AOI22X2 fu_ALU_fu_arch_U292 ( .A0(n2190), .A1(n2145), .B0(n2191), .B1(
        fu_ALU_fu_arch_N632), .Y(fu_ALU_fu_arch_n530) );
  AOI2BB2X2 U408 ( .B0(n2241), .B1(n286), .A0N(rf_RF_reg_0__12_), .A1N(n2241), 
        .Y(n837) );
  NAND2X2 U1137 ( .A(n600), .B(rf_BOOL_reg_0__0_), .Y(n599) );
  OAI211X2 fu_ALU_fu_arch_U324 ( .A0(fu_ALU_fu_arch_n462), .A1(
        fu_ALU_fu_arch_n235), .B0(fu_ALU_fu_arch_n569), .C0(
        fu_ALU_fu_arch_n570), .Y(fu_ALU_fu_arch_n567) );
  AOI2BB2X2 U404 ( .B0(n2245), .B1(n286), .A0N(fu_LSU_o1shadow_reg_12_), .A1N(
        n2246), .Y(n834) );
  OAI211X2 fu_ALU_fu_arch_U354 ( .A0(fu_ALU_fu_arch_n536), .A1(
        fu_ALU_fu_arch_n292), .B0(fu_ALU_fu_arch_n594), .C0(
        fu_ALU_fu_arch_n595), .Y(ic_socket_ALU_o1_data0_wire[17]) );
  AOI22X2 fu_ALU_fu_arch_U273 ( .A0(n2190), .A1(n2143), .B0(n2193), .B1(
        fu_ALU_fu_arch_N54), .Y(fu_ALU_fu_arch_n512) );
  CLKNAND2X8 U350 ( .A(n255), .B(n256), .Y(rf_RF_t1data_wire[15]) );
  AOI2BB2X2 U410 ( .B0(n2233), .B1(n286), .A0N(rf_RF_reg_2__12_), .A1N(n2233), 
        .Y(n839) );
  AOI22X2 U329 ( .A0(n2257), .A1(ic_socket_ALU_o1_data0_wire[16]), .B0(n2222), 
        .B1(rf_RF_reg_4__16_), .Y(n243) );
  AOI2BB2X2 U412 ( .B0(n2225), .B1(n286), .A0N(rf_RF_reg_4__12_), .A1N(n2225), 
        .Y(n841) );
  AOI2BB2X2 U438 ( .B0(n2236), .B1(n297), .A0N(rf_RF_reg_1__11_), .A1N(n2237), 
        .Y(n853) );
  AOI22X2 U406 ( .A0(n1285), .A1(n286), .B0(n283), .B1(n2244), .Y(n836) );
  AOI22X2 U435 ( .A0(n1285), .A1(n297), .B0(n294), .B1(n2244), .Y(n851) );
  AOI2BB2X2 U409 ( .B0(n2237), .B1(n286), .A0N(rf_RF_reg_1__12_), .A1N(n2237), 
        .Y(n838) );
  AOI2BB2X2 U437 ( .B0(n2240), .B1(n297), .A0N(rf_RF_reg_0__11_), .A1N(n2241), 
        .Y(n852) );
  AOI2BB2X2 U440 ( .B0(n2228), .B1(n297), .A0N(rf_RF_reg_3__11_), .A1N(n2229), 
        .Y(n855) );
  AOI2BB2X2 U439 ( .B0(n2232), .B1(n297), .A0N(rf_RF_reg_2__11_), .A1N(n2233), 
        .Y(n854) );
  AOI2BB2X2 U411 ( .B0(n2229), .B1(n286), .A0N(rf_RF_reg_3__12_), .A1N(n2229), 
        .Y(n840) );
  AOI2BB2X2 U441 ( .B0(n2224), .B1(n297), .A0N(rf_RF_reg_4__11_), .A1N(n2225), 
        .Y(n856) );
  AOI22X2 U483 ( .A0(n252), .A1(n319), .B0(fu_LSU_data_out[9]), .B1(n2248), 
        .Y(n318) );
  AOI22X2 U359 ( .A0(n252), .A1(n38), .B0(fu_LSU_data_out[14]), .B1(n2248), 
        .Y(n262) );
  AOI22X2 U367 ( .A0(n252), .A1(n65), .B0(fu_LSU_data_out[13]), .B1(n2248), 
        .Y(n270) );
  AOI22X2 U396 ( .A0(n252), .A1(n78), .B0(fu_LSU_data_out[12]), .B1(n2248), 
        .Y(n285) );
  AOI22X2 U377 ( .A0(n1285), .A1(n272), .B0(n268), .B1(n2244), .Y(n821) );
  AOI22X2 U425 ( .A0(n252), .A1(n90), .B0(fu_LSU_data_out[11]), .B1(n2248), 
        .Y(n296) );
  AOI22X2 U304 ( .A0(n2257), .A1(ic_socket_ALU_o1_data0_wire[17]), .B0(n2222), 
        .B1(rf_RF_reg_4__17_), .Y(n223) );
  AOI22X2 U454 ( .A0(fu_LSU_data_out[10]), .A1(n2248), .B0(n252), .B1(n102), 
        .Y(n307) );
  AOI2BB2X2 U382 ( .B0(n2227), .B1(n272), .A0N(rf_RF_reg_3__13_), .A1N(n2229), 
        .Y(n825) );
  AOI22X2 U337 ( .A0(n252), .A1(n30), .B0(fu_LSU_data_out[15]), .B1(n2248), 
        .Y(n251) );
  OAI211X2 fu_ALU_fu_arch_U289 ( .A0(fu_ALU_fu_arch_n388), .A1(
        fu_ALU_fu_arch_n228), .B0(fu_ALU_fu_arch_n530), .C0(
        fu_ALU_fu_arch_n531), .Y(fu_ALU_fu_arch_n525) );
  AOI2BB2X2 U383 ( .B0(n2223), .B1(n272), .A0N(rf_RF_reg_4__13_), .A1N(n2225), 
        .Y(n826) );
  AOI2BB2X2 U380 ( .B0(n2235), .B1(n272), .A0N(rf_RF_reg_1__13_), .A1N(n2237), 
        .Y(n823) );
  AOI2BB2X2 U381 ( .B0(n2231), .B1(n272), .A0N(rf_RF_reg_2__13_), .A1N(n2233), 
        .Y(n824) );
  AOI22X2 fu_ALU_fu_arch_U271 ( .A0(n2192), .A1(fu_ALU_fu_arch_N633), .B0(
        n2143), .B1(fu_ALU_fu_arch_n514), .Y(fu_ALU_fu_arch_n513) );
  AOI2BB2X2 U379 ( .B0(n2239), .B1(n272), .A0N(rf_RF_reg_0__13_), .A1N(n2241), 
        .Y(n822) );
  AOI2BB2X2 U375 ( .B0(n2245), .B1(n272), .A0N(fu_LSU_o1shadow_reg_13_), .A1N(
        n39), .Y(n819) );
  OAI211X2 fu_ALU_fu_arch_U336 ( .A0(fu_ALU_fu_arch_n316), .A1(
        fu_ALU_fu_arch_n292), .B0(fu_ALU_fu_arch_n577), .C0(
        fu_ALU_fu_arch_n578), .Y(ic_socket_ALU_o1_data0_wire[18]) );
  AOI22X2 fu_ALU_fu_arch_U257 ( .A0(n2190), .A1(n2141), .B0(n2193), .B1(
        fu_ALU_fu_arch_N55), .Y(fu_ALU_fu_arch_n495) );
  AOI2BB2X2 U346 ( .B0(n2233), .B1(n254), .A0N(rf_RF_reg_2__15_), .A1N(n2233), 
        .Y(n807) );
  AOI22X2 fu_ALU_fu_arch_U240 ( .A0(n2190), .A1(n2139), .B0(n2193), .B1(
        fu_ALU_fu_arch_N56), .Y(fu_ALU_fu_arch_n476) );
  AOI2BB2X2 U347 ( .B0(n2229), .B1(n254), .A0N(rf_RF_reg_3__15_), .A1N(n2229), 
        .Y(n808) );
  AOI22X2 U282 ( .A0(n2257), .A1(ic_socket_ALU_o1_data0_wire[18]), .B0(n2222), 
        .B1(rf_RF_reg_4__18_), .Y(n210) );
  AOI22X2 fu_ALU_fu_arch_U255 ( .A0(n2192), .A1(fu_ALU_fu_arch_N634), .B0(
        n2141), .B1(fu_ALU_fu_arch_n497), .Y(fu_ALU_fu_arch_n496) );
  AOI2BB2X2 U345 ( .B0(n2237), .B1(n254), .A0N(rf_RF_reg_1__15_), .A1N(n2237), 
        .Y(n806) );
  AOI2BB2X2 U348 ( .B0(n2225), .B1(n254), .A0N(rf_RF_reg_4__15_), .A1N(n2225), 
        .Y(n809) );
  OAI211X2 fu_ALU_fu_arch_U270 ( .A0(fu_ALU_fu_arch_n204), .A1(
        fu_ALU_fu_arch_n388), .B0(fu_ALU_fu_arch_n512), .C0(
        fu_ALU_fu_arch_n513), .Y(fu_ALU_fu_arch_n508) );
  AOI2BB2X2 U344 ( .B0(n2241), .B1(n254), .A0N(rf_RF_reg_0__15_), .A1N(n2241), 
        .Y(n805) );
  AOI2BB2X2 U341 ( .B0(n2245), .B1(n254), .A0N(fu_LSU_o1shadow_reg_15_), .A1N(
        n39), .Y(n803) );
  AOI22X2 U342 ( .A0(n1761), .A1(n254), .B0(n248), .B1(n2244), .Y(n804) );
  AOI2BB2X2 U319 ( .B0(n2245), .B1(n241), .A0N(fu_LSU_o1shadow_reg_16_), .A1N(
        n2246), .Y(n793) );
  AOI22X2 U916 ( .A0(n1761), .A1(n263), .B0(n260), .B1(n2243), .Y(n1084) );
  AOI2BB2X2 U326 ( .B0(n2224), .B1(n241), .A0N(rf_RF_reg_4__16_), .A1N(n2224), 
        .Y(n799) );
  AOI2BB2X2 U914 ( .B0(n2245), .B1(n263), .A0N(fu_LSU_o1shadow_reg_14_), .A1N(
        n39), .Y(n1082) );
  AOI22X2 fu_ALU_fu_arch_U238 ( .A0(n2191), .A1(fu_ALU_fu_arch_N635), .B0(
        n2139), .B1(fu_ALU_fu_arch_n478), .Y(fu_ALU_fu_arch_n477) );
  AOI2BB2X2 U918 ( .B0(n2239), .B1(n263), .A0N(rf_RF_reg_0__14_), .A1N(n2242), 
        .Y(n1085) );
  AOI22X2 U320 ( .A0(n1761), .A1(n241), .B0(n228), .B1(n2244), .Y(n794) );
  AOI22X2 fu_ALU_fu_arch_U222 ( .A0(n2190), .A1(n2137), .B0(n2193), .B1(
        fu_ALU_fu_arch_N57), .Y(fu_ALU_fu_arch_n453) );
  OAI211X2 fu_ALU_fu_arch_U254 ( .A0(fu_ALU_fu_arch_n187), .A1(
        fu_ALU_fu_arch_n388), .B0(fu_ALU_fu_arch_n495), .C0(
        fu_ALU_fu_arch_n496), .Y(fu_ALU_fu_arch_n489) );
  AOI2BB2X2 U920 ( .B0(n2231), .B1(n263), .A0N(rf_RF_reg_2__14_), .A1N(n2234), 
        .Y(n1087) );
  AOI2BB2X2 U919 ( .B0(n2235), .B1(n263), .A0N(rf_RF_reg_1__14_), .A1N(n2238), 
        .Y(n1086) );
  OAI211X2 U313 ( .A0(n235), .A1(n25), .B0(n236), .C0(n237), .Y(n234) );
  AOI2BB2X2 U325 ( .B0(n2228), .B1(n241), .A0N(rf_RF_reg_3__16_), .A1N(n2228), 
        .Y(n798) );
  AOI2BB2X2 U324 ( .B0(n2232), .B1(n241), .A0N(rf_RF_reg_2__16_), .A1N(n2232), 
        .Y(n797) );
  AOI2BB2X2 U921 ( .B0(n2227), .B1(n263), .A0N(rf_RF_reg_3__14_), .A1N(n2230), 
        .Y(n1088) );
  AOI22X2 U260 ( .A0(n2257), .A1(ic_socket_ALU_o1_data0_wire[19]), .B0(n2222), 
        .B1(rf_RF_reg_4__19_), .Y(n196) );
  AOI2BB2X2 U322 ( .B0(n2240), .B1(n241), .A0N(rf_RF_reg_0__16_), .A1N(n2240), 
        .Y(n795) );
  AOI2BB2X2 U922 ( .B0(n2223), .B1(n263), .A0N(rf_RF_reg_4__14_), .A1N(n2226), 
        .Y(n1089) );
  AOI2BB2X2 U323 ( .B0(n2236), .B1(n241), .A0N(rf_RF_reg_1__16_), .A1N(n2236), 
        .Y(n796) );
  AOI2BB2X2 U301 ( .B0(n2223), .B1(n221), .A0N(rf_RF_reg_4__17_), .A1N(n2224), 
        .Y(n789) );
  AOI22X2 fu_ALU_fu_arch_U205 ( .A0(n2190), .A1(n2135), .B0(n2193), .B1(
        fu_ALU_fu_arch_N58), .Y(fu_ALU_fu_arch_n431) );
  AOI32X2 U758 ( .A0(n1268), .A1(n2110), .A2(n319), .B0(n416), .B1(n2110), .Y(
        n415) );
  NAND2X2 U289 ( .A(n217), .B(n218), .Y(n781) );
  AOI22X2 U295 ( .A0(n1761), .A1(n221), .B0(n215), .B1(n2244), .Y(n784) );
  AOI2BB2X2 U300 ( .B0(n2227), .B1(n221), .A0N(rf_RF_reg_3__17_), .A1N(n2228), 
        .Y(n788) );
  AOI2BB2X2 U299 ( .B0(n2231), .B1(n221), .A0N(rf_RF_reg_2__17_), .A1N(n2232), 
        .Y(n787) );
  AOI2BB2X2 U294 ( .B0(n2245), .B1(n221), .A0N(fu_LSU_o1shadow_reg_17_), .A1N(
        n39), .Y(n783) );
  AOI22X2 fu_ALU_fu_arch_U220 ( .A0(n2191), .A1(fu_ALU_fu_arch_N636), .B0(
        n2137), .B1(fu_ALU_fu_arch_n455), .Y(fu_ALU_fu_arch_n454) );
  CLKNAND2X8 U259 ( .A(n195), .B(n196), .Y(rf_RF_t1data_wire[19]) );
  AOI2BB2X2 U297 ( .B0(n2239), .B1(n221), .A0N(rf_RF_reg_0__17_), .A1N(n2240), 
        .Y(n785) );
  AOI2BB2X2 U298 ( .B0(n2235), .B1(n221), .A0N(rf_RF_reg_1__17_), .A1N(n2236), 
        .Y(n786) );
  AOI22X2 U239 ( .A0(n2257), .A1(ic_socket_ALU_o1_data0_wire[20]), .B0(n2222), 
        .B1(rf_RF_reg_4__20_), .Y(n184) );
  AOI32X2 U747 ( .A0(n132), .A1(n411), .A2(n231), .B0(n412), .B1(n411), .Y(
        n1029) );
  AOI2BB2X2 U278 ( .B0(n2227), .B1(n208), .A0N(rf_RF_reg_3__18_), .A1N(n2229), 
        .Y(n778) );
  OAI211X2 U267 ( .A0(n203), .A1(n142), .B0(n204), .C0(n205), .Y(n771) );
  AOI2BB2X2 U277 ( .B0(n2231), .B1(n208), .A0N(rf_RF_reg_2__18_), .A1N(n2233), 
        .Y(n777) );
  AOI22X2 U273 ( .A0(n1761), .A1(n208), .B0(n201), .B1(n2243), .Y(n774) );
  INVX6 U258 ( .A(rf_RF_t1data_wire[19]), .Y(n194) );
  AOI2BB2X2 U275 ( .B0(n2239), .B1(n208), .A0N(rf_RF_reg_0__18_), .A1N(n2241), 
        .Y(n775) );
  AOI2BB2X2 U272 ( .B0(n2245), .B1(n208), .A0N(fu_LSU_o1shadow_reg_18_), .A1N(
        n39), .Y(n773) );
  NAND2X2 U757 ( .A(n414), .B(n415), .Y(n1030) );
  OAI211X2 fu_ALU_fu_arch_U219 ( .A0(fu_ALU_fu_arch_n147), .A1(
        fu_ALU_fu_arch_n430), .B0(fu_ALU_fu_arch_n453), .C0(
        fu_ALU_fu_arch_n454), .Y(fu_ALU_fu_arch_n447) );
  AOI22X2 U218 ( .A0(n2257), .A1(ic_socket_ALU_o1_data0_wire[21]), .B0(n2222), 
        .B1(rf_RF_reg_4__21_), .Y(n172) );
  AOI2BB2X2 U276 ( .B0(n2235), .B1(n208), .A0N(rf_RF_reg_1__18_), .A1N(n2237), 
        .Y(n776) );
  AOI22X2 fu_ALU_fu_arch_U203 ( .A0(n2191), .A1(fu_ALU_fu_arch_N637), .B0(
        n2135), .B1(fu_ALU_fu_arch_n433), .Y(fu_ALU_fu_arch_n432) );
  AOI2BB2X2 U279 ( .B0(n2223), .B1(n208), .A0N(rf_RF_reg_4__18_), .A1N(n2225), 
        .Y(n779) );
  AOI2BB2X2 U253 ( .B0(n2240), .B1(n194), .A0N(rf_RF_reg_0__19_), .A1N(n2240), 
        .Y(n765) );
  AOI22X2 U197 ( .A0(ic_socket_ALU_o1_bus_cntrl_wire_0_), .A1(
        ic_socket_ALU_o1_data0_wire[22]), .B0(n2222), .B1(rf_RF_reg_4__22_), 
        .Y(n160) );
  OAI2BB2X2 U675 ( .B0(n203), .B1(n1284), .A0N(fu_LSU_data_out[2]), .A1N(n2248), .Y(n979) );
  OAI2BB2X2 U648 ( .B0(n1284), .B1(n191), .A0N(fu_LSU_data_out[3]), .A1N(n2248), .Y(n964) );
  OAI2BB2X2 U621 ( .B0(n1284), .B1(n179), .A0N(fu_LSU_data_out[4]), .A1N(n2248), .Y(n949) );
  OAI2BB2X2 U567 ( .B0(n1284), .B1(n155), .A0N(fu_LSU_data_out[6]), .A1N(n2248), .Y(n919) );
  AOI2BB2X2 U255 ( .B0(n2232), .B1(n194), .A0N(rf_RF_reg_2__19_), .A1N(n2232), 
        .Y(n767) );
  OAI211X2 U246 ( .A0(n191), .A1(n142), .B0(n192), .C0(n193), .Y(n761) );
  AOI2BB2X2 U250 ( .B0(n2245), .B1(n194), .A0N(fu_LSU_o1shadow_reg_19_), .A1N(
        n39), .Y(n763) );
  OAI211X2 fu_ALU_fu_arch_U202 ( .A0(fu_ALU_fu_arch_n117), .A1(
        fu_ALU_fu_arch_n430), .B0(fu_ALU_fu_arch_n431), .C0(
        fu_ALU_fu_arch_n432), .Y(fu_ALU_fu_arch_n423) );
  OAI2BB2X2 U594 ( .B0(n1284), .B1(n167), .A0N(fu_LSU_data_out[5]), .A1N(n2248), .Y(n934) );
  AOI2BB2X2 U254 ( .B0(n2236), .B1(n194), .A0N(rf_RF_reg_1__19_), .A1N(n2236), 
        .Y(n766) );
  OAI2BB2X2 U540 ( .B0(n1284), .B1(n141), .A0N(fu_LSU_data_out[7]), .A1N(n2248), .Y(n904) );
  AOI2BB2X2 U256 ( .B0(n2228), .B1(n194), .A0N(rf_RF_reg_3__19_), .A1N(n2228), 
        .Y(n768) );
  INVX6 U237 ( .A(rf_RF_t1data_wire[20]), .Y(n182) );
  AOI2BB2X2 U257 ( .B0(n2224), .B1(n194), .A0N(rf_RF_reg_4__19_), .A1N(n2224), 
        .Y(n769) );
  AOI22X2 U251 ( .A0(n1761), .A1(n194), .B0(n189), .B1(n2243), .Y(n764) );
  AOI32X2 fu_ALU_fu_arch_U190 ( .A0(n2133), .A1(n1763), .A2(n1762), .B0(
        fu_ALU_fu_arch_N638), .B1(n2192), .Y(fu_ALU_fu_arch_n414) );
  AOI22X2 U230 ( .A0(n1761), .A1(n182), .B0(n177), .B1(n2243), .Y(n754) );
  AOI2BB2X2 U233 ( .B0(n2238), .B1(n182), .A0N(rf_RF_reg_1__20_), .A1N(n2236), 
        .Y(n756) );
  AOI2BB2X2 U236 ( .B0(n2226), .B1(n182), .A0N(rf_RF_reg_4__20_), .A1N(n2224), 
        .Y(n759) );
  AOI32X2 fu_ALU_fu_arch_U177 ( .A0(n2131), .A1(n1764), .A2(n1762), .B0(
        fu_ALU_fu_arch_N639), .B1(n2191), .Y(fu_ALU_fu_arch_n397) );
  OAI211X2 U225 ( .A0(n179), .A1(n142), .B0(n180), .C0(n181), .Y(n751) );
  AOI2BB2X2 U235 ( .B0(n2230), .B1(n182), .A0N(rf_RF_reg_3__20_), .A1N(n2228), 
        .Y(n758) );
  AOI2BB2X2 U232 ( .B0(n2242), .B1(n182), .A0N(rf_RF_reg_0__20_), .A1N(n2240), 
        .Y(n755) );
  AOI2BB2X2 U234 ( .B0(n2234), .B1(n182), .A0N(rf_RF_reg_2__20_), .A1N(n2232), 
        .Y(n757) );
  AOI22X2 U176 ( .A0(n2257), .A1(ic_socket_ALU_o1_data0_wire[23]), .B0(n2222), 
        .B1(rf_RF_reg_4__23_), .Y(n147) );
  INVX6 U216 ( .A(rf_RF_t1data_wire[21]), .Y(n170) );
  AOI2BB2X2 U229 ( .B0(n2245), .B1(n182), .A0N(fu_LSU_o1shadow_reg_20_), .A1N(
        n39), .Y(n753) );
  OAI211X2 fu_ALU_fu_arch_U210 ( .A0(fu_ALU_fu_arch_n139), .A1(
        fu_ALU_fu_arch_n388), .B0(fu_ALU_fu_arch_n442), .C0(
        fu_ALU_fu_arch_n443), .Y(ic_socket_ALU_o1_data0_wire[24]) );
  AOI22X2 fu_ALU_fu_arch_U160 ( .A0(n2190), .A1(n2130), .B0(n2191), .B1(
        fu_ALU_fu_arch_N640), .Y(fu_ALU_fu_arch_n373) );
  INVX6 U195 ( .A(rf_RF_t1data_wire[22]), .Y(n158) );
  NAND2X2 U1122 ( .A(n590), .B(n573), .Y(n588) );
  OAI211X2 U204 ( .A0(n167), .A1(n142), .B0(n168), .C0(n169), .Y(n741) );
  AOI22X2 U209 ( .A0(n1761), .A1(n170), .B0(n165), .B1(n2243), .Y(n744) );
  OAI211X2 U999 ( .A0(n536), .A1(n542), .B0(n543), .C0(n544), .Y(n541) );
  AOI2BB2X2 U208 ( .B0(n2245), .B1(n170), .A0N(fu_LSU_o1shadow_reg_21_), .A1N(
        n39), .Y(n743) );
  AOI2BB2X2 U214 ( .B0(n2229), .B1(n170), .A0N(rf_RF_reg_3__21_), .A1N(n2229), 
        .Y(n748) );
  AOI2BB2X2 U212 ( .B0(n2237), .B1(n170), .A0N(rf_RF_reg_1__21_), .A1N(n2237), 
        .Y(n746) );
  AOI2BB2X2 U215 ( .B0(n2225), .B1(n170), .A0N(rf_RF_reg_4__21_), .A1N(n2225), 
        .Y(n749) );
  AOI2BB2X2 U211 ( .B0(n2241), .B1(n170), .A0N(rf_RF_reg_0__21_), .A1N(n2241), 
        .Y(n745) );
  AOI2BB2X2 U213 ( .B0(n2233), .B1(n170), .A0N(rf_RF_reg_2__21_), .A1N(n2233), 
        .Y(n747) );
  AOI22X2 fu_ALU_fu_arch_U114 ( .A0(n2193), .A1(fu_ALU_fu_arch_N63), .B0(n2126), .B1(fu_ALU_fu_arch_n301), .Y(fu_ALU_fu_arch_n300) );
  AOI2BB2X2 U193 ( .B0(n2228), .B1(n158), .A0N(rf_RF_reg_3__22_), .A1N(n2228), 
        .Y(n738) );
  AOI2BB2X2 U192 ( .B0(n2232), .B1(n158), .A0N(rf_RF_reg_2__22_), .A1N(n2232), 
        .Y(n737) );
  AOI2BB2X2 U194 ( .B0(n2224), .B1(n158), .A0N(rf_RF_reg_4__22_), .A1N(n2224), 
        .Y(n739) );
  AOI2BB2X2 U190 ( .B0(n2240), .B1(n158), .A0N(rf_RF_reg_0__22_), .A1N(n2240), 
        .Y(n735) );
  OAI211X2 U183 ( .A0(n155), .A1(n142), .B0(n156), .C0(n157), .Y(n731) );
  AOI22X2 U188 ( .A0(n1761), .A1(n158), .B0(n153), .B1(n2243), .Y(n734) );
  INVX6 U174 ( .A(rf_RF_t1data_wire[23]), .Y(n145) );
  AOI2BB2X2 U187 ( .B0(n2245), .B1(n158), .A0N(fu_LSU_o1shadow_reg_22_), .A1N(
        n2246), .Y(n733) );
  AOI22X2 fu_ALU_fu_arch_U147 ( .A0(n2190), .A1(n2128), .B0(n2191), .B1(
        fu_ALU_fu_arch_N641), .Y(fu_ALU_fu_arch_n353) );
  AOI2BB2X2 U191 ( .B0(n2236), .B1(n158), .A0N(rf_RF_reg_1__22_), .A1N(n2236), 
        .Y(n736) );
  AO22X2 U1047 ( .A0(n1857), .A1(n553), .B0(fu_LIFTING_in1_load_wire), .B1(
        n2211), .Y(n1142) );
  INVX2 U1127 ( .A(n592), .Y(n1189) );
  OAI2BB2X2 U1121 ( .B0(n588), .B1(n578), .A0N(n2257), .A1N(n2211), .Y(n1187)
         );
  AOI2BB2X2 U169 ( .B0(n2242), .B1(n145), .A0N(rf_RF_reg_0__23_), .A1N(n2241), 
        .Y(n725) );
  AOI2BB2X2 U170 ( .B0(n2238), .B1(n145), .A0N(rf_RF_reg_1__23_), .A1N(n2237), 
        .Y(n726) );
  AOI2BB2X2 U173 ( .B0(n2226), .B1(n145), .A0N(rf_RF_reg_4__23_), .A1N(n2225), 
        .Y(n729) );
  AOI22X2 fu_ALU_fu_arch_U116 ( .A0(n2190), .A1(n2126), .B0(n2191), .B1(
        fu_ALU_fu_arch_N642), .Y(fu_ALU_fu_arch_n299) );
  AOI2BB2X2 U1084 ( .B0(n2207), .B1(n577), .A0N(ic_simm_B1_wire[1]), .A1N(
        n2207), .Y(n1163) );
  AO22X2 U1119 ( .A0(n2211), .A1(ic_socket_bool_o1_bus_cntrl_wire_0_), .B0(
        n1893), .B1(inst_decoder_instructionword_wire[35]), .Y(n1186) );
  NAND2X4 U1114 ( .A(n578), .B(n1893), .Y(n583) );
  AOI22X2 U167 ( .A0(n1761), .A1(n145), .B0(n139), .B1(n2243), .Y(n724) );
  AOI2BB2X2 U166 ( .B0(n39), .B1(n145), .A0N(fu_LSU_o1shadow_reg_23_), .A1N(
        n2246), .Y(n723) );
  AOI2BB2X2 U171 ( .B0(n2234), .B1(n145), .A0N(rf_RF_reg_2__23_), .A1N(n2233), 
        .Y(n727) );
  INVX6 U151 ( .A(rf_RF_t1data_wire[24]), .Y(n133) );
  AOI2BB2X2 U172 ( .B0(n2230), .B1(n145), .A0N(rf_RF_reg_3__23_), .A1N(n2229), 
        .Y(n728) );
  OAI211X2 U162 ( .A0(n141), .A1(n142), .B0(n143), .C0(n144), .Y(n721) );
  AOI2BB2X2 U146 ( .B0(n2240), .B1(n133), .A0N(rf_RF_reg_0__24_), .A1N(n2241), 
        .Y(n715) );
  AOI2BB2X2 U993 ( .B0(n2112), .B1(n540), .A0N(fu_ALU_t1opcode_wire[3]), .A1N(
        n2112), .Y(n1120) );
  AOI2BB2X2 U150 ( .B0(n2224), .B1(n133), .A0N(rf_RF_reg_4__24_), .A1N(n2225), 
        .Y(n719) );
  AOI2BB2X2 U149 ( .B0(n2228), .B1(n133), .A0N(rf_RF_reg_3__24_), .A1N(n2229), 
        .Y(n718) );
  AOI2BB2X2 U991 ( .B0(n2112), .B1(n531), .A0N(fu_ALU_t1opcode_wire[1]), .A1N(
        n2112), .Y(n1118) );
  AOI22X2 U1067 ( .A0(n2207), .A1(n573), .B0(n49), .B1(n2206), .Y(n1147) );
  AOI2BB2X2 U989 ( .B0(n2112), .B1(n536), .A0N(fu_ALU_t1opcode_wire[0]), .A1N(
        n2112), .Y(n1116) );
  AOI22X2 U977 ( .A0(n530), .A1(n1752), .B0(n1751), .B1(n532), .Y(n1109) );
  OAI211X2 U136 ( .A0(n125), .A1(n103), .B0(n126), .C0(n127), .Y(n711) );
  AOI2BB2X2 U987 ( .B0(n2112), .B1(n537), .A0N(fu_ALU_t1opcode_wire[2]), .A1N(
        n2112), .Y(n1114) );
  AOI22X2 U979 ( .A0(n530), .A1(n537), .B0(n527), .B1(n532), .Y(n1110) );
  AOI22X2 U1011 ( .A0(n549), .A1(n531), .B0(n547), .B1(n550), .Y(n1128) );
  AOI22X2 U1013 ( .A0(n549), .A1(n1752), .B0(n546), .B1(n550), .Y(n1129) );
  AOI2BB2X2 U147 ( .B0(n2236), .B1(n133), .A0N(rf_RF_reg_1__24_), .A1N(n2237), 
        .Y(n716) );
  INVX6 U127 ( .A(rf_RF_t1data_wire[25]), .Y(n117) );
  AOI2BB2X2 U148 ( .B0(n2232), .B1(n133), .A0N(rf_RF_reg_2__24_), .A1N(n2233), 
        .Y(n717) );
  AOI2BB2X2 U143 ( .B0(n2245), .B1(n133), .A0N(fu_LSU_o1shadow_reg_24_), .A1N(
        n2246), .Y(n713) );
  AO21X2 U997 ( .A0(fu_ALU_t1load_wire), .A1(n2211), .B0(n2112), .Y(n1122) );
  AOI22X2 U966 ( .A0(n530), .A1(n531), .B0(n239), .B1(n532), .Y(n1104) );
  AOI22X2 U144 ( .A0(n1761), .A1(n133), .B0(n123), .B1(n2243), .Y(n714) );
  AOI2BB2X2 U119 ( .B0(n39), .B1(n117), .A0N(fu_LSU_o1shadow_reg_25_), .A1N(
        n2246), .Y(n703) );
  AOI22X2 U1107 ( .A0(n581), .A1(n577), .B0(n582), .B1(n583), .Y(n1180) );
  AOI2BB2X2 U123 ( .B0(n2236), .B1(n117), .A0N(rf_RF_reg_1__25_), .A1N(n2237), 
        .Y(n706) );
  AOI22X2 U1109 ( .A0(n581), .A1(n576), .B0(n584), .B1(n583), .Y(n1181) );
  AOI2BB2X2 U126 ( .B0(n2224), .B1(n117), .A0N(rf_RF_reg_4__25_), .A1N(n2225), 
        .Y(n709) );
  AOI2BB2X2 U124 ( .B0(n2232), .B1(n117), .A0N(rf_RF_reg_2__25_), .A1N(n2233), 
        .Y(n707) );
  AOI2BB2X2 U122 ( .B0(n2240), .B1(n117), .A0N(rf_RF_reg_0__25_), .A1N(n2241), 
        .Y(n705) );
  AOI2BB2X2 U125 ( .B0(n2228), .B1(n117), .A0N(rf_RF_reg_3__25_), .A1N(n2229), 
        .Y(n708) );
  AOI22X2 U1110 ( .A0(n581), .A1(n575), .B0(n585), .B1(n583), .Y(n1182) );
  INVX6 U105 ( .A(rf_RF_t1data_wire[26]), .Y(n104) );
  AOI22X2 U120 ( .A0(n1761), .A1(n117), .B0(n110), .B1(n2243), .Y(n704) );
  AOI2BB2X2 U103 ( .B0(n2228), .B1(n104), .A0N(rf_RF_reg_3__26_), .A1N(n2230), 
        .Y(n698) );
  AOI2BB2X2 U97 ( .B0(n39), .B1(n104), .A0N(fu_LSU_o1shadow_reg_26_), .A1N(
        n2246), .Y(n693) );
  INVX6 U83 ( .A(rf_RF_t1data_wire[27]), .Y(n91) );
  AOI2BB2X2 U104 ( .B0(n2224), .B1(n104), .A0N(rf_RF_reg_4__26_), .A1N(n2226), 
        .Y(n699) );
  AOI2BB2X2 U100 ( .B0(n2240), .B1(n104), .A0N(rf_RF_reg_0__26_), .A1N(n2242), 
        .Y(n695) );
  AOI2BB2X2 U101 ( .B0(n2236), .B1(n104), .A0N(rf_RF_reg_1__26_), .A1N(n2238), 
        .Y(n696) );
  AOI22X2 U98 ( .A0(n1761), .A1(n104), .B0(n97), .B1(n2243), .Y(n694) );
  OAI211X2 fu_ALU_fu_arch_U111 ( .A0(fu_ALU_fu_arch_n291), .A1(
        fu_ALU_fu_arch_n292), .B0(fu_ALU_fu_arch_n293), .C0(
        fu_ALU_fu_arch_n294), .Y(ic_socket_ALU_o1_data0_wire[30]) );
  OAI211X2 U92 ( .A0(n99), .A1(n25), .B0(n100), .C0(n101), .Y(n691) );
  AOI2BB2X2 U102 ( .B0(n2232), .B1(n104), .A0N(rf_RF_reg_2__26_), .A1N(n2234), 
        .Y(n697) );
  AOI22X2 U76 ( .A0(n1761), .A1(n91), .B0(n85), .B1(n2243), .Y(n684) );
  OAI211X2 U71 ( .A0(n87), .A1(n25), .B0(n88), .C0(n89), .Y(n681) );
  INVX6 U62 ( .A(rf_RF_t1data_wire[28]), .Y(n79) );
  AOI2BB2X2 U75 ( .B0(n2245), .B1(n91), .A0N(fu_LSU_o1shadow_reg_27_), .A1N(
        n2245), .Y(n683) );
  AOI22X2 U49 ( .A0(fu_ALU_o1reg[28]), .A1(n2252), .B0(n2250), .B1(
        rf_RF_t1data_wire[28]), .Y(n74) );
  AOI2BB2X2 U78 ( .B0(n2240), .B1(n91), .A0N(rf_RF_reg_0__27_), .A1N(n2242), 
        .Y(n685) );
  AOI2BB2X2 U80 ( .B0(n2232), .B1(n91), .A0N(rf_RF_reg_2__27_), .A1N(n2234), 
        .Y(n687) );
  AOI2BB2X2 U82 ( .B0(n2224), .B1(n91), .A0N(rf_RF_reg_4__27_), .A1N(n2226), 
        .Y(n689) );
  AOI2BB2X2 U81 ( .B0(n2228), .B1(n91), .A0N(rf_RF_reg_3__27_), .A1N(n2230), 
        .Y(n688) );
  AOI2BB2X2 U79 ( .B0(n2236), .B1(n91), .A0N(rf_RF_reg_1__27_), .A1N(n2238), 
        .Y(n686) );
  AOI2BB2X2 U58 ( .B0(n2236), .B1(n79), .A0N(rf_RF_reg_1__28_), .A1N(n2238), 
        .Y(n676) );
  AOI2BB2X2 U54 ( .B0(n39), .B1(n79), .A0N(fu_LSU_o1shadow_reg_28_), .A1N(n39), 
        .Y(n673) );
  AOI2BB2X2 U59 ( .B0(n2232), .B1(n79), .A0N(rf_RF_reg_2__28_), .A1N(n2234), 
        .Y(n677) );
  AOI2BB2X2 U60 ( .B0(n2228), .B1(n79), .A0N(rf_RF_reg_3__28_), .A1N(n2230), 
        .Y(n678) );
  AOI2BB2X2 U57 ( .B0(n2240), .B1(n79), .A0N(rf_RF_reg_0__28_), .A1N(n2242), 
        .Y(n675) );
  OAI211X2 U50 ( .A0(n75), .A1(n25), .B0(n76), .C0(n77), .Y(n671) );
  AOI22X2 U55 ( .A0(n1761), .A1(n79), .B0(n73), .B1(n2243), .Y(n674) );
  AOI2BB2X2 U61 ( .B0(n2224), .B1(n79), .A0N(rf_RF_reg_4__28_), .A1N(n2226), 
        .Y(n679) );
  AOI22X2 U30 ( .A0(n2123), .A1(n1861), .B0(n29), .B1(n65), .Y(n64) );
  INVX6 U41 ( .A(n1861), .Y(n66) );
  AOI22X2 U28 ( .A0(fu_ALU_o1reg[29]), .A1(n2252), .B0(n2250), .B1(n1861), .Y(
        n61) );
  INVX6 U20 ( .A(n1862), .Y(n40) );
  INVX6 U939 ( .A(n1860), .Y(n512) );
  AOI22X2 U2 ( .A0(fu_ALU_o1reg[31]), .A1(n2252), .B0(n2250), .B1(n1860), .Y(
        n21) );
  AOI22X2 U34 ( .A0(n1761), .A1(n66), .B0(n60), .B1(n2243), .Y(n664) );
  AOI22X2 U4 ( .A0(n2123), .A1(n1860), .B0(n29), .B1(n30), .Y(n27) );
  AOI2BB2X2 U39 ( .B0(n2228), .B1(n66), .A0N(rf_RF_reg_3__29_), .A1N(n2230), 
        .Y(n668) );
  OAI211X2 U29 ( .A0(n62), .A1(n25), .B0(n63), .C0(n64), .Y(n661) );
  AOI2BB2X2 U38 ( .B0(n2232), .B1(n66), .A0N(rf_RF_reg_2__29_), .A1N(n2234), 
        .Y(n667) );
  AOI2BB2X2 U37 ( .B0(n2236), .B1(n66), .A0N(rf_RF_reg_1__29_), .A1N(n2238), 
        .Y(n666) );
  AOI2BB2X2 U40 ( .B0(n2224), .B1(n66), .A0N(rf_RF_reg_4__29_), .A1N(n2226), 
        .Y(n669) );
  AOI2BB2X2 U33 ( .B0(n39), .B1(n66), .A0N(fu_LSU_o1shadow_reg_29_), .A1N(n39), 
        .Y(n663) );
  AOI22X2 U9 ( .A0(n2123), .A1(n1862), .B0(n29), .B1(n38), .Y(n37) );
  AOI22X2 U7 ( .A0(fu_ALU_fu_arch_sub_200_B_30_), .A1(n2252), .B0(n2250), .B1(
        n1862), .Y(n34) );
  AOI2BB2X2 U36 ( .B0(n2240), .B1(n66), .A0N(rf_RF_reg_0__29_), .A1N(n2242), 
        .Y(n665) );
  AOI2BB2X2 U15 ( .B0(n2240), .B1(n40), .A0N(rf_RF_reg_0__30_), .A1N(n2239), 
        .Y(n655) );
  AOI2BB2X2 U937 ( .B0(n2227), .B1(n512), .A0N(rf_RF_reg_3__31_), .A1N(n2230), 
        .Y(n1096) );
  AOI2BB2X2 U18 ( .B0(n2228), .B1(n40), .A0N(rf_RF_reg_3__30_), .A1N(n2227), 
        .Y(n658) );
  AOI2BB2X2 U12 ( .B0(n39), .B1(n40), .A0N(fu_LSU_o1shadow_reg_30_), .A1N(
        n2245), .Y(n653) );
  AOI2BB2X2 U17 ( .B0(n2232), .B1(n40), .A0N(rf_RF_reg_2__30_), .A1N(n2231), 
        .Y(n657) );
  AOI2BB2X2 U935 ( .B0(n2235), .B1(n512), .A0N(rf_RF_reg_1__31_), .A1N(n2238), 
        .Y(n1094) );
  AOI2BB2X2 U934 ( .B0(n2239), .B1(n512), .A0N(rf_RF_reg_0__31_), .A1N(n2242), 
        .Y(n1093) );
  AOI2BB2X2 U19 ( .B0(n2224), .B1(n40), .A0N(rf_RF_reg_4__30_), .A1N(n2223), 
        .Y(n659) );
  AOI2BB2X2 U936 ( .B0(n2231), .B1(n512), .A0N(rf_RF_reg_2__31_), .A1N(n2234), 
        .Y(n1095) );
  AOI2BB2X2 U931 ( .B0(n2245), .B1(n512), .A0N(fu_LSU_o1shadow_reg_31_), .A1N(
        n2246), .Y(n1091) );
  AOI2BB2X2 U16 ( .B0(n2236), .B1(n40), .A0N(rf_RF_reg_1__30_), .A1N(n2235), 
        .Y(n656) );
  OAI211X2 U3 ( .A0(n24), .A1(n25), .B0(n26), .C0(n27), .Y(n649) );
  AOI2BB2X2 U938 ( .B0(n2223), .B1(n512), .A0N(rf_RF_reg_4__31_), .A1N(n2226), 
        .Y(n1097) );
  AOI22X2 U932 ( .A0(n1761), .A1(n512), .B0(n20), .B1(n2244), .Y(n1092) );
  AOI22X2 U13 ( .A0(n1761), .A1(n40), .B0(n33), .B1(n2243), .Y(n654) );
  OAI211X2 U8 ( .A0(n35), .A1(n25), .B0(n36), .C0(n37), .Y(n651) );
  AOI22X2 U926 ( .A0(n1777), .A1(rf_RF_reg_2__14_), .B0(n2218), .B1(
        rf_RF_reg_3__14_), .Y(n509) );
  AOI22X2 U1152 ( .A0(n1777), .A1(rf_RF_reg_2__0_), .B0(n2219), .B1(
        rf_RF_reg_0__0_), .Y(n610) );
  AOI22X2 U642 ( .A0(n1777), .A1(rf_RF_reg_2__4_), .B0(n2218), .B1(
        rf_RF_reg_3__4_), .Y(n380) );
  AOI222X2 U111 ( .A0(ic_socket_lsu_o1_data0_wire[26]), .A1(n2187), .B0(n1777), 
        .B1(rf_RF_reg_2__26_), .C0(n2256), .C1(
        ic_socket_LIFTING_o1_data0_wire[26]), .Y(n108) );
  AOI22X2 U1271 ( .A0(n1777), .A1(rf_RF_reg_2__1_), .B0(n2218), .B1(
        rf_RF_reg_3__1_), .Y(n629) );
  AOI22X2 U669 ( .A0(n1777), .A1(rf_RF_reg_2__3_), .B0(n2218), .B1(
        rf_RF_reg_3__3_), .Y(n390) );
  AOI22X2 U615 ( .A0(n1777), .A1(rf_RF_reg_2__5_), .B0(n2218), .B1(
        rf_RF_reg_3__5_), .Y(n370) );
  AOI22X2 U698 ( .A0(n1777), .A1(rf_RF_reg_2__2_), .B0(n2218), .B1(
        rf_RF_reg_3__2_), .Y(n400) );
  AOI22X2 U943 ( .A0(n1777), .A1(rf_RF_reg_2__31_), .B0(n2256), .B1(
        ic_socket_LIFTING_o1_data0_wire[31]), .Y(n518) );
  AOI222X2 U89 ( .A0(ic_socket_lsu_o1_data0_wire[27]), .A1(n2187), .B0(n1777), 
        .B1(rf_RF_reg_2__27_), .C0(n2256), .C1(
        ic_socket_LIFTING_o1_data0_wire[27]), .Y(n95) );
  CLKNAND2X2 fu_ALU_fu_arch_U564 ( .A(n2162), .B(n2188), .Y(
        fu_ALU_fu_arch_n726) );
  CLKNAND2X2 fu_ALU_fu_arch_U520 ( .A(n2160), .B(n2188), .Y(
        fu_ALU_fu_arch_n704) );
  AOI32X2 fu_ALU_fu_arch_U345 ( .A0(n2149), .A1(n2148), .A2(n1762), .B0(n2190), 
        .B1(n2149), .Y(fu_ALU_fu_arch_n586) );
  CLKNAND2X2 fu_ALU_fu_arch_U144 ( .A(n2197), .B(fu_ALU_o1reg[29]), .Y(
        fu_ALU_fu_arch_n349) );
  NAND2X2 fu_ALU_fu_arch_U598 ( .A(n2202), .B(n1780), .Y(fu_ALU_fu_arch_n371)
         );
  CLKNAND2X2 fu_ALU_fu_arch_U584 ( .A(n2197), .B(fu_ALU_fu_arch_sub_200_B_14_), 
        .Y(fu_ALU_fu_arch_n731) );
  NAND2X5 fu_ALU_fu_arch_U651 ( .A(fu_ALU_fu_arch_n249), .B(
        fu_ALU_fu_arch_n612), .Y(fu_ALU_fu_arch_n235) );
  AOI22X2 fu_ALU_fu_arch_U544 ( .A0(n2198), .A1(n2138), .B0(n2201), .B1(n1780), 
        .Y(fu_ALU_fu_arch_n713) );
  CLKNAND2X2 fu_ALU_fu_arch_U536 ( .A(n2200), .B(n2151), .Y(
        fu_ALU_fu_arch_n710) );
  CLKNAND2X2 fu_ALU_fu_arch_U523 ( .A(n2200), .B(n2157), .Y(
        fu_ALU_fu_arch_n706) );
  AOI22X2 fu_ALU_fu_arch_U196 ( .A0(n2197), .A1(n1780), .B0(n2200), .B1(
        fu_ALU_o1reg[24]), .Y(fu_ALU_fu_arch_n421) );
  INVX4 fu_ALU_fu_arch_U484 ( .A(n2103), .Y(fu_ALU_fu_arch_n136) );
  AOI22X2 fu_ALU_fu_arch_U208 ( .A0(n1775), .A1(fu_ALU_fu_arch_n438), .B0(
        fu_ALU_fu_arch_n249), .B1(fu_ALU_fu_arch_n435), .Y(fu_ALU_fu_arch_n436) );
  AOI22X2 fu_ALU_fu_arch_U427 ( .A0(n1775), .A1(n1888), .B0(
        fu_ALU_fu_arch_n249), .B1(n1842), .Y(fu_ALU_fu_arch_n652) );
  AOI22X2 fu_ALU_fu_arch_U407 ( .A0(n1775), .A1(n1830), .B0(
        fu_ALU_fu_arch_n249), .B1(n1841), .Y(fu_ALU_fu_arch_n637) );
  AOI22X2 fu_ALU_fu_arch_U442 ( .A0(n1775), .A1(n1837), .B0(
        fu_ALU_fu_arch_n249), .B1(n1845), .Y(fu_ALU_fu_arch_n665) );
  AOI222X2 fu_ALU_fu_arch_U155 ( .A0(fu_ALU_fu_arch_n366), .A1(n1775), .B0(
        n1840), .B1(n2105), .C0(n1795), .C1(n2104), .Y(fu_ALU_fu_arch_n365) );
  INVX2 fu_ALU_fu_arch_U333 ( .A(fu_ALU_fu_arch_n574), .Y(fu_ALU_fu_arch_n575)
         );
  AOI222X2 fu_ALU_fu_arch_U123 ( .A0(fu_ALU_fu_arch_n313), .A1(n1775), .B0(
        n1794), .B1(n2104), .C0(n1801), .C1(n2105), .Y(fu_ALU_fu_arch_n306) );
  OAI21X1 fu_ALU_fu_arch_U134 ( .A0(fu_ALU_fu_arch_n331), .A1(
        fu_ALU_fu_arch_sub_200_B_not_2_), .B0(fu_ALU_fu_arch_n332), .Y(
        fu_ALU_fu_arch_n330) );
  AOI222X2 fu_ALU_fu_arch_U142 ( .A0(fu_ALU_fu_arch_n345), .A1(n1775), .B0(
        n1796), .B1(n2105), .C0(n1882), .C1(n2104), .Y(fu_ALU_fu_arch_n344) );
  OAI2B11X2 fu_ALU_fu_arch_U73 ( .A1N(fu_ALU_fu_arch_n214), .A0(
        fu_ALU_fu_arch_n212), .B0(fu_ALU_fu_arch_n215), .C0(
        fu_ALU_fu_arch_n216), .Y(ic_socket_ALU_o1_data0_wire[4]) );
  OAI211X2 fu_ALU_fu_arch_U124 ( .A0(fu_ALU_fu_arch_n316), .A1(
        fu_ALU_fu_arch_n212), .B0(fu_ALU_fu_arch_n317), .C0(
        fu_ALU_fu_arch_n318), .Y(ic_socket_ALU_o1_data0_wire[2]) );
  AOI221X2 U590 ( .A0(n2186), .A1(ic_socket_gcu_o1_data0_wire[6]), .B0(n2257), 
        .B1(ic_socket_ALU_o1_data0_wire[6]), .C0(n362), .Y(n358) );
  AOI221X2 U563 ( .A0(n2186), .A1(ic_socket_gcu_o1_data0_wire[7]), .B0(n2257), 
        .B1(ic_socket_ALU_o1_data0_wire[7]), .C0(n352), .Y(n348) );
  AOI221X2 U507 ( .A0(n2186), .A1(ic_socket_gcu_o1_data0_wire[9]), .B0(n2257), 
        .B1(ic_socket_ALU_o1_data0_wire[9]), .C0(n328), .Y(n324) );
  AOI221X2 fu_ALU_fu_arch_U502 ( .A0(n2160), .A1(fu_ALU_fu_arch_n153), .B0(
        fu_ALU_fu_arch_n696), .B1(fu_ALU_o1reg[11]), .C0(fu_ALU_fu_arch_n697), 
        .Y(fu_ALU_fu_arch_n695) );
  AOI221X2 U478 ( .A0(n2186), .A1(ic_socket_gcu_o1_data0_wire[10]), .B0(n2257), 
        .B1(ic_socket_ALU_o1_data0_wire[10]), .C0(n315), .Y(n311) );
  NAND4X2 fu_ALU_fu_arch_U501 ( .A(fu_ALU_fu_arch_n692), .B(
        fu_ALU_fu_arch_n693), .C(fu_ALU_fu_arch_n694), .D(fu_ALU_fu_arch_n695), 
        .Y(ic_socket_ALU_o1_data0_wire[11]) );
  AOI221X2 U420 ( .A0(n2186), .A1(ic_socket_gcu_o1_data0_wire[12]), .B0(n2257), 
        .B1(ic_socket_ALU_o1_data0_wire[12]), .C0(n293), .Y(n289) );
  NAND2X2 fu_ALU_fu_arch_U383 ( .A(fu_ALU_fu_arch_n615), .B(
        fu_ALU_fu_arch_n616), .Y(fu_ALU_fu_arch_n614) );
  AOI221X2 U391 ( .A0(n2186), .A1(ic_socket_gcu_o1_data0_wire[13]), .B0(n2257), 
        .B1(ic_socket_ALU_o1_data0_wire[13]), .C0(n282), .Y(n278) );
  AOI22X2 U603 ( .A0(n1285), .A1(n365), .B0(n363), .B1(n2244), .Y(n941) );
  OAI22X1 U1136 ( .A0(inst_decoder_instructionword_wire[40]), .A1(n599), .B0(
        inst_decoder_instructionword_wire[39]), .B1(n600), .Y(n598) );
  OAI211X2 fu_ALU_fu_arch_U193 ( .A0(fu_ALU_fu_arch_n107), .A1(
        fu_ALU_fu_arch_n388), .B0(fu_ALU_fu_arch_n418), .C0(
        fu_ALU_fu_arch_n419), .Y(ic_socket_ALU_o1_data0_wire[25]) );
  AOI22X2 U107 ( .A0(n2257), .A1(ic_socket_ALU_o1_data0_wire[26]), .B0(n2221), 
        .B1(rf_RF_reg_4__26_), .Y(n106) );
  AOI22X2 U85 ( .A0(n2257), .A1(ic_socket_ALU_o1_data0_wire[27]), .B0(n2221), 
        .B1(rf_RF_reg_4__27_), .Y(n93) );
  OAI211X2 fu_ALU_fu_arch_U139 ( .A0(fu_ALU_fu_arch_n337), .A1(
        fu_ALU_fu_arch_n270), .B0(fu_ALU_fu_arch_n338), .C0(
        fu_ALU_fu_arch_n339), .Y(ic_socket_ALU_o1_data0_wire[29]) );
  AOI22X2 U22 ( .A0(n2257), .A1(ic_socket_ALU_o1_data0_wire[30]), .B0(n2221), 
        .B1(rf_RF_reg_4__30_), .Y(n51) );
  INVX5 fu_ALU_fu_arch_U710 ( .A(fu_ALU_opc1reg[0]), .Y(fu_ALU_fu_arch_n746)
         );
  CLKINVX24 fu_ALU_fu_arch_U655 ( .A(n2106), .Y(fu_ALU_fu_arch_n249) );
  CLKNAND2X2 U794 ( .A(ic_socket_lsu_o1_data0_wire[7]), .B(n2212), .Y(n451) );
  OAI22X1 fu_ALU_fu_arch_U19 ( .A0(fu_ALU_fu_arch_n131), .A1(
        fu_ALU_fu_arch_n132), .B0(fu_ALU_fu_arch_n133), .B1(
        fu_ALU_fu_arch_n134), .Y(fu_ALU_fu_arch_n114) );
  NOR3X2 fu_ALU_fu_arch_U436 ( .A(fu_ALU_fu_arch_n659), .B(fu_ALU_fu_arch_n660), .C(fu_ALU_fu_arch_n661), .Y(fu_ALU_fu_arch_n656) );
  AOI31X1 U1135 ( .A0(inst_decoder_instructionword_wire[40]), .A1(
        inst_decoder_instructionword_wire[39]), .A2(n597), .B0(n598), .Y(n596)
         );
  CLKNAND2X8 U238 ( .A(n183), .B(n184), .Y(rf_RF_t1data_wire[20]) );
  CLKNAND2X8 U217 ( .A(n171), .B(n172), .Y(rf_RF_t1data_wire[21]) );
  CLKNAND2X8 U196 ( .A(n159), .B(n160), .Y(rf_RF_t1data_wire[22]) );
  NAND2X2 fu_ALU_fu_arch_U188 ( .A(fu_ALU_fu_arch_n414), .B(
        fu_ALU_fu_arch_n415), .Y(fu_ALU_fu_arch_n406) );
  CLKNAND2X8 U175 ( .A(n146), .B(n147), .Y(rf_RF_t1data_wire[23]) );
  NAND2X2 fu_ALU_fu_arch_U175 ( .A(fu_ALU_fu_arch_n397), .B(
        fu_ALU_fu_arch_n398), .Y(fu_ALU_fu_arch_n385) );
  AOI22X2 U155 ( .A0(n2257), .A1(ic_socket_ALU_o1_data0_wire[24]), .B0(n2222), 
        .B1(rf_RF_reg_4__24_), .Y(n135) );
  ADDFX1 fu_ALU_fu_arch_sub_200_U2_30 ( .A(n2126), .B(
        fu_ALU_fu_arch_sub_200_B_not_30_), .CI(
        fu_ALU_fu_arch_sub_200_carry_30_), .CO(
        fu_ALU_fu_arch_sub_200_carry_31_), .S(fu_ALU_fu_arch_N642) );
  CLKNAND2X8 U152 ( .A(n134), .B(n135), .Y(rf_RF_t1data_wire[24]) );
  ADDFX1 fu_ALU_fu_arch_add_171_U1_30 ( .A(n2126), .B(
        fu_ALU_fu_arch_sub_200_B_30_), .CI(fu_ALU_fu_arch_add_171_carry_30_), 
        .CO(fu_ALU_fu_arch_add_171_carry_31_), .S(fu_ALU_fu_arch_N63) );
  AOI22X2 U129 ( .A0(n2257), .A1(ic_socket_ALU_o1_data0_wire[25]), .B0(n2221), 
        .B1(rf_RF_reg_4__25_), .Y(n119) );
  CLKNAND2X8 U128 ( .A(n118), .B(n119), .Y(rf_RF_t1data_wire[25]) );
  CLKNAND2X8 U106 ( .A(n105), .B(n106), .Y(rf_RF_t1data_wire[26]) );
  AOI22X2 U64 ( .A0(n2257), .A1(ic_socket_ALU_o1_data0_wire[28]), .B0(n2221), 
        .B1(rf_RF_reg_4__28_), .Y(n81) );
  CLKNAND2X8 U84 ( .A(n92), .B(n93), .Y(rf_RF_t1data_wire[27]) );
  AOI22X2 U43 ( .A0(n2257), .A1(ic_socket_ALU_o1_data0_wire[29]), .B0(n2221), 
        .B1(rf_RF_reg_4__29_), .Y(n69) );
  CLKNAND2X2 U1056 ( .A(inst_decoder_N121), .B(n537), .Y(n568) );
  OR2X2 fu_ALU_fu_arch_U698 ( .A(n1779), .B(fu_ALU_fu_arch_sub_200_A_1_), .Y(
        fu_ALU_fu_arch_n250) );
  AOI21X1 fu_ALU_fu_arch_U398 ( .A0(fu_ALU_o1reg[31]), .A1(fu_ALU_fu_arch_n111), .B0(fu_ALU_fu_arch_n290), .Y(fu_ALU_fu_arch_n352) );
  INVX6 fu_ALU_fu_arch_U652 ( .A(fu_ALU_fu_arch_n108), .Y(fu_ALU_fu_arch_n612)
         );
  INVX5 fu_ALU_fu_arch_U607 ( .A(fu_ALU_fu_arch_n208), .Y(fu_ALU_fu_arch_n169)
         );
  OAI22X1 fu_ALU_fu_arch_U72 ( .A0(fu_ALU_fu_arch_n133), .A1(
        fu_ALU_fu_arch_n132), .B0(fu_ALU_fu_arch_n137), .B1(
        fu_ALU_fu_arch_n134), .Y(fu_ALU_fu_arch_n200) );
  AOI211X2 fu_ALU_fu_arch_U332 ( .A0(n2104), .A1(fu_ALU_fu_arch_n481), .B0(
        fu_ALU_fu_arch_n518), .C0(fu_ALU_fu_arch_n575), .Y(fu_ALU_fu_arch_n262) );
  AOI21X2 fu_ALU_fu_arch_U300 ( .A0(fu_ALU_fu_arch_n178), .A1(
        fu_ALU_fu_arch_n539), .B0(fu_ALU_fu_arch_n540), .Y(fu_ALU_fu_arch_n538) );
  AOI221X2 U644 ( .A0(n2186), .A1(ic_socket_gcu_o1_data0_wire[4]), .B0(n2257), 
        .B1(ic_socket_ALU_o1_data0_wire[4]), .C0(n382), .Y(n378) );
  ADDFX2 fu_ALU_fu_arch_add_171_U1_21 ( .A(n2143), .B(
        fu_ALU_fu_arch_sub_200_B_21_), .CI(fu_ALU_fu_arch_add_171_carry_21_), 
        .CO(fu_ALU_fu_arch_add_171_carry_22_), .S(fu_ALU_fu_arch_N54) );
  ADDFX1 fu_ALU_fu_arch_add_171_U1_26 ( .A(n2133), .B(n2132), .CI(
        fu_ALU_fu_arch_add_171_carry_26_), .CO(
        fu_ALU_fu_arch_add_171_carry_27_), .S(fu_ALU_fu_arch_N59) );
  ADDFX1 fu_ALU_fu_arch_add_171_U1_27 ( .A(n2131), .B(
        fu_ALU_fu_arch_sub_200_B_27_), .CI(fu_ALU_fu_arch_add_171_carry_27_), 
        .CO(fu_ALU_fu_arch_add_171_carry_28_), .S(fu_ALU_fu_arch_N60) );
  ADDFX1 fu_ALU_fu_arch_add_171_U1_28 ( .A(n2130), .B(
        fu_ALU_fu_arch_lt_gt_188_A_28_), .CI(fu_ALU_fu_arch_add_171_carry_28_), 
        .CO(fu_ALU_fu_arch_add_171_carry_29_), .S(fu_ALU_fu_arch_N61) );
  CLKNAND2X8 U63 ( .A(n80), .B(n81), .Y(rf_RF_t1data_wire[28]) );
  CLKNAND2X2 fu_ALU_fu_arch_U470 ( .A(n2202), .B(n2151), .Y(
        fu_ALU_fu_arch_n674) );
  AOI21X1 fu_ALU_fu_arch_U301 ( .A0(fu_ALU_fu_arch_n292), .A1(
        fu_ALU_fu_arch_n430), .B0(fu_ALU_fu_arch_n541), .Y(fu_ALU_fu_arch_n540) );
  ADDFX1 fu_ALU_fu_arch_add_171_U1_24 ( .A(n2137), .B(fu_ALU_o1reg[24]), .CI(
        fu_ALU_fu_arch_add_171_carry_24_), .CO(
        fu_ALU_fu_arch_add_171_carry_25_), .S(fu_ALU_fu_arch_N57) );
  ADDFX1 fu_ALU_fu_arch_add_171_U1_25 ( .A(n2135), .B(fu_ALU_o1reg[25]), .CI(
        fu_ALU_fu_arch_add_171_carry_25_), .CO(
        fu_ALU_fu_arch_add_171_carry_26_), .S(fu_ALU_fu_arch_N58) );
  ADDFX1 fu_ALU_fu_arch_sub_200_U2_26 ( .A(n2133), .B(n1763), .CI(
        fu_ALU_fu_arch_sub_200_carry_26_), .CO(
        fu_ALU_fu_arch_sub_200_carry_27_), .S(fu_ALU_fu_arch_N638) );
  ADDFX1 fu_ALU_fu_arch_sub_200_U2_27 ( .A(n2131), .B(n1764), .CI(
        fu_ALU_fu_arch_sub_200_carry_27_), .CO(
        fu_ALU_fu_arch_sub_200_carry_28_), .S(fu_ALU_fu_arch_N639) );
  DFFSRX4 inst_fetch_pc_reg_reg_1_ ( .D(n1028), .CK(clk), .SN(n1027), .RN(
        n1026), .Q(inst_fetch_pc_reg_1_), .QN(n1295) );
  DFFSRX4 inst_fetch_pc_reg_reg_4_ ( .D(n952), .CK(clk), .SN(n951), .RN(n950), 
        .Q(inst_fetch_pc_reg_4_), .QN(n1301) );
  DFFSRX4 inst_fetch_pc_reg_reg_6_ ( .D(n922), .CK(clk), .SN(n921), .RN(n920), 
        .Q(inst_fetch_pc_reg_6_), .QN(n1305) );
  DFFSRX4 inst_fetch_pc_reg_reg_2_ ( .D(n982), .CK(clk), .SN(n981), .RN(n980), 
        .Q(inst_fetch_pc_reg_2_), .QN(n1297) );
  DFFSRX4 inst_fetch_pc_reg_reg_7_ ( .D(n907), .CK(clk), .SN(n906), .RN(n905), 
        .Q(inst_fetch_pc_reg_7_), .QN(n1307) );
  DFFSRX4 inst_fetch_pc_reg_reg_3_ ( .D(n967), .CK(clk), .SN(n966), .RN(n965), 
        .Q(inst_fetch_pc_reg_3_), .QN(n1299) );
  DFFSRX4 inst_fetch_pc_reg_reg_0_ ( .D(n1077), .CK(clk), .SN(n1076), .RN(
        n1075), .Q(inst_fetch_pc_reg_0_), .QN(inst_fetch_increased_pc_0_) );
  DFFSRX4 inst_fetch_pc_reg_reg_8_ ( .D(n892), .CK(clk), .SN(n891), .RN(n890), 
        .Q(inst_fetch_pc_reg_8_), .QN(n1293) );
  DFFSRX4 inst_fetch_pc_reg_reg_5_ ( .D(n937), .CK(clk), .SN(n936), .RN(n935), 
        .Q(inst_fetch_pc_reg_5_), .QN(n1303) );
  DFFSRX4 inst_fetch_pc_reg_reg_9_ ( .D(n877), .CK(clk), .SN(n876), .RN(n875), 
        .Q(inst_fetch_pc_reg_9_), .QN(n1309) );
  DFFSRX4 inst_fetch_pc_reg_reg_10_ ( .D(n862), .CK(clk), .SN(n861), .RN(n860), 
        .Q(inst_fetch_pc_reg_10_), .QN(n1311) );
  DFFSRX4 inst_fetch_pc_reg_reg_12_ ( .D(n832), .CK(clk), .SN(n831), .RN(n830), 
        .Q(inst_fetch_pc_reg_12_), .QN(n1315) );
  DFFSRX4 inst_fetch_pc_reg_reg_11_ ( .D(n847), .CK(clk), .SN(n846), .RN(n845), 
        .Q(inst_fetch_pc_reg_11_), .QN(n1313) );
  DFFSRX4 inst_fetch_pc_reg_reg_13_ ( .D(n817), .CK(clk), .SN(n816), .RN(n815), 
        .Q(inst_fetch_pc_reg_13_), .QN(n1317) );
  DFFSRX4 inst_fetch_pc_reg_reg_14_ ( .D(n1080), .CK(clk), .SN(n1079), .RN(
        n1078), .Q(inst_fetch_pc_reg_14_), .QN(n1319) );
  DFFRX4 inst_fetch_instruction_reg_reg_6_ ( .D(n1227), .CK(clk), .RN(rstx), 
        .Q(inst_decoder_instructionword_wire[6]), .QN(n576) );
  DFFRX4 inst_fetch_instruction_reg_reg_0_ ( .D(n1233), .CK(clk), .RN(rstx), 
        .Q(inst_decoder_N119), .QN(n536) );
  DFFRX4 fu_LSU_status_addr_reg_reg_1__0_ ( .D(n1102), .CK(clk), .RN(rstx), 
        .Q(fu_LSU_status_addr_reg_1__0_), .QN(n454) );
  DFFRX4 fu_ALU_o1reg_reg_1_ ( .D(n993), .CK(clk), .RN(rstx), .Q(
        fu_ALU_o1reg[1]), .QN(n1738) );
  DFFRX4 fu_ALU_o1reg_reg_2_ ( .D(n978), .CK(clk), .RN(rstx), .Q(
        fu_ALU_o1reg[2]), .QN(n2175) );
  DFFRX4 fu_ALU_t1reg_reg_0_ ( .D(n1121), .CK(clk), .RN(rstx), .QN(n2184) );
  DFFRX4 fu_LSU_o1shadow_reg_reg_9_ ( .D(n879), .CK(clk), .RN(rstx), .Q(
        fu_LSU_o1shadow_reg_9_) );
  DFFRX4 fu_ALU_t1reg_reg_13_ ( .D(n818), .CK(clk), .RN(rstx), .Q(
        fu_ALU_t1reg[13]), .QN(n1740) );
  DFFRX4 fu_ALU_o1reg_reg_18_ ( .D(n770), .CK(clk), .RN(rstx), .QN(n2148) );
  DFFRX4 fu_ALU_t1reg_reg_21_ ( .D(n742), .CK(clk), .RN(rstx), .Q(
        fu_ALU_t1reg[21]), .QN(n1736) );
  DFFRX4 inst_decoder_fu_ALU_in2_load_reg_reg ( .D(n1144), .CK(clk), .RN(rstx), 
        .QN(n521) );
  DFFRX4 inst_decoder_fu_LIFTING_x1_load_reg_reg ( .D(n1142), .CK(clk), .RN(
        rstx), .Q(fu_LIFTING_in1_load_wire), .QN(n1757) );
  DFFRX4 fu_ALU_t1reg_reg_23_ ( .D(n722), .CK(clk), .RN(rstx), .Q(
        fu_ALU_t1reg[23]), .QN(n1737) );
  DFFRX4 inst_decoder_fu_LSU_in1t_load_reg_reg ( .D(n1112), .CK(clk), .RN(rstx), .Q(fu_LSU_t1load_wire), .QN(n524) );
  DFFRX4 inst_decoder_fu_LSU_opc_reg_reg_0_ ( .D(n1109), .CK(clk), .RN(rstx), 
        .QN(n2182) );
  DFFRX4 fu_ALU_t1reg_reg_31_ ( .D(n1090), .CK(clk), .RN(rstx), .Q(
        fu_ALU_t1reg[31]), .QN(n1739) );
  DFFRX4 fu_ALU_o1reg_reg_30_ ( .D(n650), .CK(clk), .RN(rstx), .QN(n2125) );
  DFFRX2 inst_fetch_instruction_reg_reg_5_ ( .D(n1228), .CK(clk), .RN(rstx), 
        .Q(inst_decoder_instructionword_wire[5]), .QN(n551) );
  DFFRX2 inst_decoder_simm_cntrl_B1_reg_reg_0_ ( .D(n1179), .CK(clk), .RN(rstx), .Q(ic_simm_cntrl_B1_wire_0_), .QN(n2259) );
  DFFRX2 inst_decoder_socket_RF_o1_bus_cntrl_reg_reg_0_ ( .D(n1183), .CK(clk), 
        .RN(rstx), .Q(ic_socket_RF_o1_bus_cntrl_wire_0_), .QN(n586) );
  DFFRQX2 fu_ALU_o1reg_reg_26_ ( .D(n690), .CK(clk), .RN(rstx), .Q(
        fu_ALU_o1reg[26]) );
  DFFRQX4 fu_ALU_o1reg_reg_28_ ( .D(n670), .CK(clk), .RN(rstx), .Q(
        fu_ALU_o1reg[28]) );
  DFFRX2 fu_ALU_t1reg_reg_28_ ( .D(n672), .CK(clk), .RN(rstx), .Q(
        fu_ALU_t1reg[28]), .QN(n1747) );
  DFFRX1 fu_ALU_o1reg_reg_15_ ( .D(n800), .CK(clk), .RN(rstx), .Q(
        fu_ALU_o1reg[15]), .QN(n1746) );
  DFFRX2 fu_ALU_t1reg_reg_9_ ( .D(n878), .CK(clk), .RN(rstx), .Q(
        fu_ALU_t1reg[9]), .QN(n1745) );
  DFFRX2 fu_ALU_t1reg_reg_12_ ( .D(n833), .CK(clk), .RN(rstx), .Q(
        fu_ALU_t1reg[12]), .QN(n1744) );
  DFFRX1 fu_ALU_o1reg_reg_7_ ( .D(n903), .CK(clk), .RN(rstx), .Q(
        fu_ALU_o1reg[7]), .QN(n1743) );
  DFFRX2 fu_ALU_t1reg_reg_8_ ( .D(n893), .CK(clk), .RN(rstx), .Q(
        fu_ALU_t1reg[8]), .QN(n1742) );
  DFFRX2 fu_ALU_t1reg_reg_6_ ( .D(n923), .CK(clk), .RN(rstx), .Q(
        fu_ALU_t1reg[6]), .QN(n1741) );
  DFFRQX4 fu_LSU_status_addr_reg_reg_1__1_ ( .D(n1065), .CK(clk), .RN(rstx), 
        .Q(fu_LSU_status_addr_reg_1__1_) );
  DFFRQX2 fu_LSU_o1shadow_reg_reg_15_ ( .D(n803), .CK(clk), .RN(rstx), .Q(
        fu_LSU_o1shadow_reg_15_) );
  DFFRQX4 fu_ALU_o1reg_reg_4_ ( .D(n948), .CK(clk), .RN(rstx), .Q(
        fu_ALU_o1reg[4]) );
  DFFRQX4 fu_ALU_o1reg_reg_19_ ( .D(n760), .CK(clk), .RN(rstx), .Q(
        fu_ALU_o1reg[19]) );
  DFFRQX4 fu_ALU_o1reg_reg_8_ ( .D(n888), .CK(clk), .RN(rstx), .Q(
        fu_ALU_o1reg[8]) );
  DFFRQX4 inst_fetch_reset_cntr_reg_0_ ( .D(n1248), .CK(clk), .RN(rstx), .Q(
        inst_fetch_reset_cntr_0_) );
  DFFRQX4 inst_decoder_fu_LSU_in2_load_reg_reg ( .D(n1133), .CK(clk), .RN(rstx), .Q(fu_LSU_o1load_wire) );
  DFFRQX4 inst_fetch_reset_cntr_reg_10_ ( .D(n1243), .CK(clk), .RN(rstx), .Q(
        inst_fetch_reset_cntr_10_) );
  DFFRQX2 fu_ALU_t1reg_reg_4_ ( .D(n953), .CK(clk), .RN(rstx), .Q(
        fu_ALU_t1reg[4]) );
  DFFRX2 inst_fetch_instruction_reg_reg_33_ ( .D(n1200), .CK(clk), .RN(rstx), 
        .Q(inst_decoder_instructionword_wire[33]) );
  DFFRX2 inst_fetch_instruction_reg_reg_31_ ( .D(n1202), .CK(clk), .RN(rstx), 
        .Q(inst_decoder_instructionword_wire[31]) );
  DFFRX2 inst_fetch_instruction_reg_reg_29_ ( .D(n1204), .CK(clk), .RN(rstx), 
        .Q(inst_decoder_instructionword_wire[29]) );
  DFFRX2 inst_fetch_instruction_reg_reg_25_ ( .D(n1208), .CK(clk), .RN(rstx), 
        .Q(inst_decoder_instructionword_wire[25]) );
  DFFRX2 inst_fetch_instruction_reg_reg_9_ ( .D(n1224), .CK(clk), .RN(rstx), 
        .Q(inst_decoder_instructionword_wire[9]) );
  DFFRX2 inst_fetch_instruction_reg_reg_8_ ( .D(n1225), .CK(clk), .RN(rstx), 
        .Q(inst_decoder_instructionword_wire[8]), .QN(n575) );
  DFFRX2 inst_fetch_instruction_reg_reg_7_ ( .D(n1226), .CK(clk), .RN(rstx), 
        .Q(inst_decoder_instructionword_wire[7]), .QN(n577) );
  DFFRX2 inst_fetch_instruction_reg_reg_34_ ( .D(n1199), .CK(clk), .RN(rstx), 
        .Q(inst_decoder_instructionword_wire[34]) );
  DFFRX2 inst_fetch_instruction_reg_reg_32_ ( .D(n1201), .CK(clk), .RN(rstx), 
        .Q(inst_decoder_instructionword_wire[32]) );
  DFFRX2 inst_fetch_instruction_reg_reg_30_ ( .D(n1203), .CK(clk), .RN(rstx), 
        .Q(inst_decoder_instructionword_wire[30]) );
  DFFRX2 inst_fetch_instruction_reg_reg_28_ ( .D(n1205), .CK(clk), .RN(rstx), 
        .Q(inst_decoder_instructionword_wire[28]) );
  DFFRX2 inst_fetch_instruction_reg_reg_27_ ( .D(n1206), .CK(clk), .RN(rstx), 
        .Q(inst_decoder_instructionword_wire[27]) );
  DFFRX2 inst_fetch_instruction_reg_reg_26_ ( .D(n1207), .CK(clk), .RN(rstx), 
        .Q(inst_decoder_instructionword_wire[26]) );
  DFFRX2 inst_fetch_instruction_reg_reg_24_ ( .D(n1209), .CK(clk), .RN(rstx), 
        .Q(inst_decoder_instructionword_wire[24]) );
  DFFRX2 inst_fetch_instruction_reg_reg_23_ ( .D(n1210), .CK(clk), .RN(rstx), 
        .Q(inst_decoder_instructionword_wire[23]) );
  DFFRX2 inst_fetch_instruction_reg_reg_22_ ( .D(n1211), .CK(clk), .RN(rstx), 
        .Q(inst_decoder_instructionword_wire[22]) );
  DFFRX2 inst_fetch_instruction_reg_reg_21_ ( .D(n1212), .CK(clk), .RN(rstx), 
        .Q(inst_decoder_instructionword_wire[21]) );
  DFFRX2 inst_fetch_instruction_reg_reg_20_ ( .D(n1213), .CK(clk), .RN(rstx), 
        .Q(inst_decoder_instructionword_wire[20]) );
  DFFRX2 inst_fetch_instruction_reg_reg_19_ ( .D(n1214), .CK(clk), .RN(rstx), 
        .Q(inst_decoder_instructionword_wire[19]) );
  DFFRX2 inst_fetch_instruction_reg_reg_18_ ( .D(n1215), .CK(clk), .RN(rstx), 
        .Q(inst_decoder_instructionword_wire[18]) );
  DFFRX2 inst_fetch_instruction_reg_reg_17_ ( .D(n1216), .CK(clk), .RN(rstx), 
        .Q(inst_decoder_instructionword_wire[17]) );
  DFFRX2 inst_fetch_instruction_reg_reg_16_ ( .D(n1217), .CK(clk), .RN(rstx), 
        .Q(inst_decoder_instructionword_wire[16]) );
  DFFRX2 inst_fetch_instruction_reg_reg_15_ ( .D(n1218), .CK(clk), .RN(rstx), 
        .Q(inst_decoder_instructionword_wire[15]) );
  DFFRX2 inst_fetch_instruction_reg_reg_14_ ( .D(n1219), .CK(clk), .RN(rstx), 
        .Q(inst_decoder_instructionword_wire[14]) );
  DFFRX2 inst_fetch_instruction_reg_reg_13_ ( .D(n1220), .CK(clk), .RN(rstx), 
        .Q(inst_decoder_instructionword_wire[13]) );
  DFFRX2 inst_fetch_instruction_reg_reg_12_ ( .D(n1221), .CK(clk), .RN(rstx), 
        .Q(inst_decoder_instructionword_wire[12]) );
  DFFRX2 inst_fetch_instruction_reg_reg_11_ ( .D(n1222), .CK(clk), .RN(rstx), 
        .Q(inst_decoder_instructionword_wire[11]) );
  DFFRX2 inst_fetch_instruction_reg_reg_10_ ( .D(n1223), .CK(clk), .RN(rstx), 
        .Q(inst_decoder_instructionword_wire[10]) );
  DFFRX1 inst_fetch_pc_prev_reg_reg_14_ ( .D(imem_addr[14]), .CK(clk), .RN(
        rstx), .QN(n1318) );
  DFFRX1 inst_fetch_pc_prev_reg_reg_13_ ( .D(imem_addr[13]), .CK(clk), .RN(
        rstx), .QN(n1316) );
  DFFRX1 inst_fetch_pc_prev_reg_reg_12_ ( .D(imem_addr[12]), .CK(clk), .RN(
        rstx), .QN(n1314) );
  DFFRX1 inst_fetch_pc_prev_reg_reg_11_ ( .D(imem_addr[11]), .CK(clk), .RN(
        rstx), .QN(n1312) );
  DFFRX1 inst_fetch_pc_prev_reg_reg_10_ ( .D(imem_addr[10]), .CK(clk), .RN(
        rstx), .QN(n1310) );
  DFFRX1 inst_fetch_pc_prev_reg_reg_9_ ( .D(imem_addr[9]), .CK(clk), .RN(rstx), 
        .QN(n1308) );
  DFFRX1 inst_fetch_pc_prev_reg_reg_7_ ( .D(imem_addr[7]), .CK(clk), .RN(rstx), 
        .QN(n1306) );
  DFFRX1 inst_fetch_pc_prev_reg_reg_6_ ( .D(imem_addr[6]), .CK(clk), .RN(rstx), 
        .QN(n1304) );
  DFFRX1 inst_fetch_pc_prev_reg_reg_5_ ( .D(imem_addr[5]), .CK(clk), .RN(rstx), 
        .QN(n1302) );
  DFFRX1 inst_fetch_pc_prev_reg_reg_4_ ( .D(imem_addr[4]), .CK(clk), .RN(rstx), 
        .QN(n1300) );
  DFFRX1 inst_fetch_pc_prev_reg_reg_3_ ( .D(imem_addr[3]), .CK(clk), .RN(rstx), 
        .QN(n1298) );
  DFFRX1 inst_fetch_pc_prev_reg_reg_2_ ( .D(imem_addr[2]), .CK(clk), .RN(rstx), 
        .QN(n1296) );
  DFFRX1 inst_fetch_pc_prev_reg_reg_1_ ( .D(imem_addr[1]), .CK(clk), .RN(rstx), 
        .QN(n1294) );
  DFFRX1 inst_fetch_pc_prev_reg_reg_8_ ( .D(imem_addr[8]), .CK(clk), .RN(rstx), 
        .QN(n1292) );
  DFFRX1 inst_fetch_pc_prev_reg_reg_0_ ( .D(imem_addr[0]), .CK(clk), .RN(rstx), 
        .QN(n1291) );
  DFFRX2 fu_LSU_status_addr_reg_reg_0__2_ ( .D(n1101), .CK(clk), .RN(rstx), 
        .Q(fu_LSU_status_addr_reg_0__2_) );
  DFFRX2 fu_LSU_status_addr_reg_reg_0__3_ ( .D(n1108), .CK(clk), .RN(rstx), 
        .QN(n535) );
  DFFRX2 fu_LSU_status_addr_reg_reg_0__4_ ( .D(n1106), .CK(clk), .RN(rstx), 
        .QN(n533) );
  DFFRX2 fu_ALU_t1reg_reg_1_ ( .D(n1031), .CK(clk), .RN(rstx), .QN(n2178) );
  DFFRX2 fu_LSU_addr_reg_reg_2_ ( .D(n955), .CK(clk), .RN(rstx), .Q(
        fu_LSU_addr[2]) );
  DFFRX2 fu_LSU_status_addr_reg_reg_0__1_ ( .D(n1066), .CK(clk), .RN(rstx), 
        .QN(n499) );
  DFFRX2 rf_RF_reg_reg_4__1_ ( .D(n1072), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_4__1_) );
  DFFRX2 rf_RF_reg_reg_3__1_ ( .D(n1071), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_3__1_) );
  DFFRX2 rf_RF_reg_reg_2__1_ ( .D(n1070), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_2__1_) );
  DFFRX2 rf_RF_reg_reg_1__1_ ( .D(n1069), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_1__1_) );
  DFFRX2 rf_RF_reg_reg_0__1_ ( .D(n1068), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_0__1_) );
  DFFRX2 fu_ALU_o1temp_reg_1_ ( .D(n1067), .CK(clk), .RN(rstx), .QN(n403) );
  DFFRX2 fu_LSU_addr_reg_reg_4_ ( .D(n925), .CK(clk), .RN(rstx), .Q(
        fu_LSU_addr[4]) );
  DFFRX2 inst_fetch_return_addr_reg_reg_1_ ( .D(n1073), .CK(clk), .RN(rstx), 
        .Q(ic_socket_gcu_o1_data0_wire[1]) );
  DFFRX2 fu_LSU_addr_reg_reg_0_ ( .D(n985), .CK(clk), .RN(rstx), .Q(
        fu_LSU_addr[0]) );
  DFFRX1 fu_ALU_t1reg_reg_2_ ( .D(n983), .CK(clk), .RN(rstx), .Q(
        fu_ALU_t1reg[2]) );
  DFFRX2 fu_LSU_r1_reg_reg_14_ ( .D(n1047), .CK(clk), .RN(rstx), .Q(
        ic_socket_lsu_o1_data0_wire[14]) );
  DFFRX2 fu_LSU_r1_reg_reg_13_ ( .D(n1046), .CK(clk), .RN(rstx), .Q(
        ic_socket_lsu_o1_data0_wire[13]) );
  DFFRX2 fu_LSU_r1_reg_reg_12_ ( .D(n1045), .CK(clk), .RN(rstx), .Q(
        ic_socket_lsu_o1_data0_wire[12]) );
  DFFRX2 fu_LSU_r1_reg_reg_11_ ( .D(n1044), .CK(clk), .RN(rstx), .Q(
        ic_socket_lsu_o1_data0_wire[11]) );
  DFFRX2 fu_LSU_r1_reg_reg_10_ ( .D(n1043), .CK(clk), .RN(rstx), .Q(
        ic_socket_lsu_o1_data0_wire[10]) );
  DFFRX2 fu_LSU_r1_reg_reg_9_ ( .D(n1042), .CK(clk), .RN(rstx), .Q(
        ic_socket_lsu_o1_data0_wire[9]) );
  DFFRX2 fu_LSU_r1_reg_reg_8_ ( .D(n1041), .CK(clk), .RN(rstx), .Q(
        ic_socket_lsu_o1_data0_wire[8]) );
  DFFRX2 fu_LSU_addr_reg_reg_5_ ( .D(n910), .CK(clk), .RN(rstx), .Q(
        fu_LSU_addr[5]) );
  DFFRX1 fu_ALU_t1reg_reg_7_ ( .D(n908), .CK(clk), .RN(rstx), .Q(
        fu_ALU_t1reg[7]) );
  DFFRX2 fu_ALU_o1temp_reg_4_ ( .D(n956), .CK(clk), .RN(rstx), .QN(n373) );
  DFFRX2 rf_RF_reg_reg_4__4_ ( .D(n961), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_4__4_) );
  DFFRX2 rf_RF_reg_reg_3__4_ ( .D(n960), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_3__4_) );
  DFFRX2 rf_RF_reg_reg_2__4_ ( .D(n959), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_2__4_) );
  DFFRX2 rf_RF_reg_reg_1__4_ ( .D(n958), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_1__4_) );
  DFFRX2 rf_RF_reg_reg_0__4_ ( .D(n957), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_0__4_) );
  DFFRX2 fu_LSU_o1shadow_reg_reg_4_ ( .D(n954), .CK(clk), .RN(rstx), .Q(
        fu_LSU_o1shadow_reg_4_) );
  DFFRX2 fu_ALU_o1temp_reg_6_ ( .D(n926), .CK(clk), .RN(rstx), .QN(n353) );
  DFFRX2 rf_RF_reg_reg_4__6_ ( .D(n931), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_4__6_) );
  DFFRX2 rf_RF_reg_reg_3__6_ ( .D(n930), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_3__6_) );
  DFFRX2 rf_RF_reg_reg_2__6_ ( .D(n929), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_2__6_) );
  DFFRX2 rf_RF_reg_reg_1__6_ ( .D(n928), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_1__6_) );
  DFFRX2 rf_RF_reg_reg_0__6_ ( .D(n927), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_0__6_) );
  DFFRX2 fu_LSU_o1shadow_reg_reg_6_ ( .D(n924), .CK(clk), .RN(rstx), .Q(
        fu_LSU_o1shadow_reg_6_) );
  DFFRX2 fu_LSU_r1_reg_reg_7_ ( .D(n1040), .CK(clk), .RN(rstx), .Q(
        ic_socket_lsu_o1_data0_wire[7]) );
  DFFRX2 fu_LSU_r1_reg_reg_6_ ( .D(n1039), .CK(clk), .RN(rstx), .Q(
        ic_socket_lsu_o1_data0_wire[6]) );
  DFFRX2 fu_LSU_r1_reg_reg_5_ ( .D(n1038), .CK(clk), .RN(rstx), .Q(
        ic_socket_lsu_o1_data0_wire[5]) );
  DFFRX2 fu_LSU_r1_reg_reg_4_ ( .D(n1037), .CK(clk), .RN(rstx), .Q(
        ic_socket_lsu_o1_data0_wire[4]) );
  DFFRX2 fu_LSU_r1_reg_reg_3_ ( .D(n1036), .CK(clk), .RN(rstx), .Q(
        ic_socket_lsu_o1_data0_wire[3]) );
  DFFRX2 fu_LSU_r1_reg_reg_2_ ( .D(n1035), .CK(clk), .RN(rstx), .Q(
        ic_socket_lsu_o1_data0_wire[2]) );
  DFFRX2 fu_LSU_r1_reg_reg_1_ ( .D(n1034), .CK(clk), .RN(rstx), .Q(
        ic_socket_lsu_o1_data0_wire[1]) );
  DFFRX2 fu_LSU_r1_reg_reg_0_ ( .D(n1033), .CK(clk), .RN(rstx), .Q(
        ic_socket_lsu_o1_data0_wire[0]) );
  DFFRX2 fu_LSU_r1_reg_reg_15_ ( .D(n1048), .CK(clk), .RN(rstx), .Q(
        ic_socket_lsu_o1_data0_wire[15]) );
  DFFRX2 inst_fetch_return_addr_reg_reg_4_ ( .D(n962), .CK(clk), .RN(rstx), 
        .Q(ic_socket_gcu_o1_data0_wire[4]) );
  DFFRX2 rf_RF_reg_reg_4__2_ ( .D(n991), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_4__2_) );
  DFFRX2 rf_RF_reg_reg_3__2_ ( .D(n990), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_3__2_) );
  DFFRX2 rf_RF_reg_reg_2__2_ ( .D(n989), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_2__2_) );
  DFFRX2 rf_RF_reg_reg_1__2_ ( .D(n988), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_1__2_) );
  DFFRX2 rf_RF_reg_reg_0__2_ ( .D(n987), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_0__2_) );
  DFFRX2 fu_ALU_o1temp_reg_2_ ( .D(n986), .CK(clk), .RN(rstx), .QN(n393) );
  DFFRX2 fu_LSU_o1shadow_reg_reg_2_ ( .D(n984), .CK(clk), .RN(rstx), .Q(
        fu_LSU_o1shadow_reg_2_) );
  DFFRX2 inst_fetch_return_addr_reg_reg_6_ ( .D(n932), .CK(clk), .RN(rstx), 
        .Q(ic_socket_gcu_o1_data0_wire[6]) );
  DFFRX2 fu_LSU_addr_reg_reg_1_ ( .D(n970), .CK(clk), .RN(rstx), .Q(
        fu_LSU_addr[1]) );
  DFFRX1 fu_ALU_t1reg_reg_3_ ( .D(n968), .CK(clk), .RN(rstx), .Q(
        fu_ALU_t1reg[3]) );
  DFFRX2 fu_ALU_o1temp_reg_7_ ( .D(n911), .CK(clk), .RN(rstx), .QN(n342) );
  DFFRX2 rf_RF_reg_reg_4__7_ ( .D(n916), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_4__7_) );
  DFFRX2 rf_RF_reg_reg_3__7_ ( .D(n915), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_3__7_) );
  DFFRX2 rf_RF_reg_reg_2__7_ ( .D(n914), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_2__7_) );
  DFFRX2 rf_RF_reg_reg_1__7_ ( .D(n913), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_1__7_) );
  DFFRX2 rf_RF_reg_reg_0__7_ ( .D(n912), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_0__7_) );
  DFFRX2 fu_LSU_o1shadow_reg_reg_7_ ( .D(n909), .CK(clk), .RN(rstx), .Q(
        fu_LSU_o1shadow_reg_7_) );
  DFFRX2 inst_fetch_return_addr_reg_reg_2_ ( .D(n992), .CK(clk), .RN(rstx), 
        .Q(ic_socket_gcu_o1_data0_wire[2]) );
  DFFRX2 inst_fetch_return_addr_reg_reg_7_ ( .D(n917), .CK(clk), .RN(rstx), 
        .Q(ic_socket_gcu_o1_data0_wire[7]) );
  DFFRX2 fu_LSU_addr_reg_reg_3_ ( .D(n940), .CK(clk), .RN(rstx), .Q(
        fu_LSU_addr[3]) );
  DFFRX2 fu_LSU_addr_reg_reg_6_ ( .D(n895), .CK(clk), .RN(rstx), .Q(
        fu_LSU_addr[6]) );
  DFFRX2 fu_LSU_r1_reg_reg_30_ ( .D(n1063), .CK(clk), .RN(rstx), .Q(
        ic_socket_lsu_o1_data0_wire[30]) );
  DFFRX2 fu_LSU_r1_reg_reg_29_ ( .D(n1062), .CK(clk), .RN(rstx), .Q(
        ic_socket_lsu_o1_data0_wire[29]) );
  DFFRX2 fu_LSU_r1_reg_reg_28_ ( .D(n1061), .CK(clk), .RN(rstx), .Q(
        ic_socket_lsu_o1_data0_wire[28]) );
  DFFRX2 fu_LSU_r1_reg_reg_27_ ( .D(n1060), .CK(clk), .RN(rstx), .Q(
        ic_socket_lsu_o1_data0_wire[27]) );
  DFFRX2 fu_LSU_r1_reg_reg_26_ ( .D(n1059), .CK(clk), .RN(rstx), .Q(
        ic_socket_lsu_o1_data0_wire[26]) );
  DFFRX2 fu_LSU_r1_reg_reg_25_ ( .D(n1058), .CK(clk), .RN(rstx), .Q(
        ic_socket_lsu_o1_data0_wire[25]) );
  DFFRX2 fu_LSU_r1_reg_reg_24_ ( .D(n1057), .CK(clk), .RN(rstx), .Q(
        ic_socket_lsu_o1_data0_wire[24]) );
  DFFRX2 fu_LSU_r1_reg_reg_31_ ( .D(n1064), .CK(clk), .RN(rstx), .QN(n491) );
  DFFRX2 fu_LSU_r1_reg_reg_23_ ( .D(n1056), .CK(clk), .RN(rstx), .QN(n150) );
  DFFRX2 fu_LSU_r1_reg_reg_22_ ( .D(n1055), .CK(clk), .RN(rstx), .QN(n162) );
  DFFRX2 fu_LSU_r1_reg_reg_21_ ( .D(n1054), .CK(clk), .RN(rstx), .QN(n174) );
  DFFRX2 fu_LSU_r1_reg_reg_20_ ( .D(n1053), .CK(clk), .RN(rstx), .QN(n186) );
  DFFRX2 fu_LSU_r1_reg_reg_19_ ( .D(n1052), .CK(clk), .RN(rstx), .QN(n198) );
  DFFRX2 fu_LSU_r1_reg_reg_18_ ( .D(n1051), .CK(clk), .RN(rstx), .QN(n212) );
  DFFRX2 fu_LSU_r1_reg_reg_17_ ( .D(n1050), .CK(clk), .RN(rstx), .QN(n225) );
  DFFRX2 fu_LSU_r1_reg_reg_16_ ( .D(n1049), .CK(clk), .RN(rstx), .QN(n245) );
  DFFRX2 rf_RF_reg_reg_4__3_ ( .D(n976), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_4__3_) );
  DFFRX2 rf_RF_reg_reg_3__3_ ( .D(n975), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_3__3_) );
  DFFRX2 rf_RF_reg_reg_2__3_ ( .D(n974), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_2__3_) );
  DFFRX2 rf_RF_reg_reg_1__3_ ( .D(n973), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_1__3_) );
  DFFRX2 rf_RF_reg_reg_0__3_ ( .D(n972), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_0__3_) );
  DFFRX2 fu_ALU_o1temp_reg_3_ ( .D(n971), .CK(clk), .RN(rstx), .QN(n383) );
  DFFRX2 fu_LSU_o1shadow_reg_reg_3_ ( .D(n969), .CK(clk), .RN(rstx), .Q(
        fu_LSU_o1shadow_reg_3_) );
  DFFRX2 rf_BOOL_reg_reg_1__0_ ( .D(n1190), .CK(clk), .RN(rstx), .Q(
        rf_BOOL_reg_1__0_), .QN(n604) );
  DFFRX2 inst_fetch_return_addr_reg_reg_3_ ( .D(n977), .CK(clk), .RN(rstx), 
        .Q(ic_socket_gcu_o1_data0_wire[3]) );
  DFFRX2 fu_LSU_addr_reg_reg_7_ ( .D(n880), .CK(clk), .RN(rstx), .Q(
        fu_LSU_addr[7]) );
  DFFRX2 fu_ALU_o1temp_reg_0_ ( .D(n1143), .CK(clk), .RN(rstx), .QN(n519) );
  DFFRX2 fu_LSU_status_addr_reg_reg_0__0_ ( .D(n1103), .CK(clk), .RN(rstx), 
        .QN(n529) );
  DFFRX1 fu_ALU_o1reg_reg_5_ ( .D(n933), .CK(clk), .RN(rstx), .Q(
        fu_ALU_o1reg[5]), .QN(n2170) );
  DFFRX2 fu_ALU_o1temp_reg_5_ ( .D(n941), .CK(clk), .RN(rstx), .QN(n363) );
  DFFRX2 rf_RF_reg_reg_4__5_ ( .D(n946), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_4__5_) );
  DFFRX2 rf_RF_reg_reg_3__5_ ( .D(n945), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_3__5_) );
  DFFRX2 rf_RF_reg_reg_2__5_ ( .D(n944), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_2__5_) );
  DFFRX2 rf_RF_reg_reg_1__5_ ( .D(n943), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_1__5_) );
  DFFRX2 rf_RF_reg_reg_0__5_ ( .D(n942), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_0__5_) );
  DFFRX2 fu_LSU_o1shadow_reg_reg_5_ ( .D(n939), .CK(clk), .RN(rstx), .Q(
        fu_LSU_o1shadow_reg_5_) );
  DFFRX2 rf_RF_reg_reg_4__0_ ( .D(n1127), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_4__0_) );
  DFFRX2 rf_RF_reg_reg_3__0_ ( .D(n1126), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_3__0_) );
  DFFRX2 rf_RF_reg_reg_2__0_ ( .D(n1125), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_2__0_) );
  DFFRX2 rf_RF_reg_reg_1__0_ ( .D(n1124), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_1__0_) );
  DFFRX2 rf_RF_reg_reg_0__0_ ( .D(n1123), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_0__0_) );
  DFFRX2 inst_fetch_return_addr_reg_reg_8_ ( .D(n902), .CK(clk), .RN(rstx), 
        .Q(ic_socket_gcu_o1_data0_wire[8]) );
  DFFRX2 inst_fetch_return_addr_reg_reg_0_ ( .D(n1074), .CK(clk), .RN(rstx), 
        .Q(ic_socket_gcu_o1_data0_wire[0]) );
  DFFRX2 inst_fetch_return_addr_reg_reg_5_ ( .D(n947), .CK(clk), .RN(rstx), 
        .Q(ic_socket_gcu_o1_data0_wire[5]) );
  DFFRX2 fu_LSU_addr_reg_reg_8_ ( .D(n865), .CK(clk), .RN(rstx), .Q(
        fu_LSU_addr[8]) );
  DFFRX1 fu_ALU_t1reg_reg_10_ ( .D(n863), .CK(clk), .RN(rstx), .Q(
        fu_ALU_t1reg[10]) );
  DFFRX2 fu_ALU_o1temp_reg_8_ ( .D(n896), .CK(clk), .RN(rstx), .QN(n329) );
  DFFRX2 rf_RF_reg_reg_4__8_ ( .D(n901), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_4__8_) );
  DFFRX2 rf_RF_reg_reg_3__8_ ( .D(n900), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_3__8_) );
  DFFRX2 rf_RF_reg_reg_2__8_ ( .D(n899), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_2__8_) );
  DFFRX2 rf_RF_reg_reg_1__8_ ( .D(n898), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_1__8_) );
  DFFRX2 rf_RF_reg_reg_0__8_ ( .D(n897), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_0__8_) );
  DFFRX2 fu_LSU_o1shadow_reg_reg_8_ ( .D(n894), .CK(clk), .RN(rstx), .Q(
        fu_LSU_o1shadow_reg_8_) );
  DFFRX1 fu_ALU_o1reg_reg_9_ ( .D(n873), .CK(clk), .RN(rstx), .Q(
        fu_ALU_o1reg[9]) );
  DFFRX2 fu_ALU_o1temp_reg_9_ ( .D(n881), .CK(clk), .RN(rstx), .QN(n316) );
  DFFRX2 rf_RF_reg_reg_4__9_ ( .D(n886), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_4__9_) );
  DFFRX2 rf_RF_reg_reg_3__9_ ( .D(n885), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_3__9_) );
  DFFRX2 rf_RF_reg_reg_2__9_ ( .D(n884), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_2__9_) );
  DFFRX2 rf_RF_reg_reg_1__9_ ( .D(n883), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_1__9_) );
  DFFRX2 rf_RF_reg_reg_0__9_ ( .D(n882), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_0__9_) );
  DFFRX2 inst_fetch_return_addr_reg_reg_9_ ( .D(n887), .CK(clk), .RN(rstx), 
        .Q(ic_socket_gcu_o1_data0_wire[9]) );
  DFFRX2 fu_LSU_addr_reg_reg_10_ ( .D(n835), .CK(clk), .RN(rstx), .Q(
        fu_LSU_addr[10]) );
  DFFRX2 fu_ALU_o1temp_reg_10_ ( .D(n866), .CK(clk), .RN(rstx), .QN(n305) );
  DFFRX2 rf_RF_reg_reg_4__10_ ( .D(n871), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_4__10_) );
  DFFRX2 rf_RF_reg_reg_3__10_ ( .D(n870), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_3__10_) );
  DFFRX2 rf_RF_reg_reg_2__10_ ( .D(n869), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_2__10_) );
  DFFRX2 rf_RF_reg_reg_1__10_ ( .D(n868), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_1__10_) );
  DFFRX2 rf_RF_reg_reg_0__10_ ( .D(n867), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_0__10_) );
  DFFRX2 fu_LSU_o1shadow_reg_reg_10_ ( .D(n864), .CK(clk), .RN(rstx), .Q(
        fu_LSU_o1shadow_reg_10_) );
  DFFRX2 fu_LSU_addr_reg_reg_9_ ( .D(n850), .CK(clk), .RN(rstx), .Q(
        fu_LSU_addr[9]) );
  DFFRX1 fu_ALU_t1reg_reg_11_ ( .D(n848), .CK(clk), .RN(rstx), .Q(
        fu_ALU_t1reg[11]) );
  DFFRX2 fu_LSU_data_out_reg_reg_8_ ( .D(n889), .CK(clk), .RN(rstx), .Q(
        fu_LSU_data_out[8]) );
  DFFRX2 inst_fetch_return_addr_reg_reg_10_ ( .D(n872), .CK(clk), .RN(rstx), 
        .Q(ic_socket_gcu_o1_data0_wire[10]) );
  DFFRX2 fu_ALU_o1temp_reg_12_ ( .D(n836), .CK(clk), .RN(rstx), .QN(n283) );
  DFFRX2 rf_RF_reg_reg_4__12_ ( .D(n841), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_4__12_) );
  DFFRX2 rf_RF_reg_reg_3__12_ ( .D(n840), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_3__12_) );
  DFFRX2 rf_RF_reg_reg_2__12_ ( .D(n839), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_2__12_) );
  DFFRX2 rf_RF_reg_reg_1__12_ ( .D(n838), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_1__12_) );
  DFFRX2 rf_RF_reg_reg_0__12_ ( .D(n837), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_0__12_) );
  DFFRX2 fu_LSU_o1shadow_reg_reg_12_ ( .D(n834), .CK(clk), .RN(rstx), .Q(
        fu_LSU_o1shadow_reg_12_) );
  DFFRX2 fu_LSU_data_out_reg_reg_1_ ( .D(n1030), .CK(clk), .RN(rstx), .Q(
        fu_LSU_data_out[1]) );
  DFFRX2 fu_LSU_data_out_reg_reg_0_ ( .D(n1029), .CK(clk), .RN(rstx), .Q(
        fu_LSU_data_out[0]) );
  DFFRX2 fu_LSU_data_out_reg_reg_12_ ( .D(n829), .CK(clk), .RN(rstx), .Q(
        fu_LSU_data_out[12]) );
  DFFRX2 fu_LSU_data_out_reg_reg_9_ ( .D(n874), .CK(clk), .RN(rstx), .Q(
        fu_LSU_data_out[9]) );
  DFFRX2 fu_LSU_data_out_reg_reg_10_ ( .D(n859), .CK(clk), .RN(rstx), .Q(
        fu_LSU_data_out[10]) );
  DFFRX2 fu_ALU_o1temp_reg_11_ ( .D(n851), .CK(clk), .RN(rstx), .QN(n294) );
  DFFRX2 rf_RF_reg_reg_4__11_ ( .D(n856), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_4__11_) );
  DFFRX2 rf_RF_reg_reg_3__11_ ( .D(n855), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_3__11_) );
  DFFRX2 rf_RF_reg_reg_2__11_ ( .D(n854), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_2__11_) );
  DFFRX2 rf_RF_reg_reg_1__11_ ( .D(n853), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_1__11_) );
  DFFRX2 rf_RF_reg_reg_0__11_ ( .D(n852), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_0__11_) );
  DFFRX2 fu_LSU_o1shadow_reg_reg_11_ ( .D(n849), .CK(clk), .RN(rstx), .Q(
        fu_LSU_o1shadow_reg_11_) );
  DFFRX2 inst_fetch_return_addr_reg_reg_12_ ( .D(n842), .CK(clk), .RN(rstx), 
        .Q(ic_socket_gcu_o1_data0_wire[12]) );
  DFFRX2 fu_LSU_data_out_reg_reg_11_ ( .D(n844), .CK(clk), .RN(rstx), .Q(
        fu_LSU_data_out[11]) );
  DFFRX1 fu_ALU_t1reg_reg_15_ ( .D(n802), .CK(clk), .RN(rstx), .Q(
        fu_ALU_t1reg[15]) );
  DFFRX2 fu_LSU_addr_reg_reg_11_ ( .D(n820), .CK(clk), .RN(rstx), .Q(
        fu_LSU_addr[11]) );
  DFFRX2 inst_fetch_return_addr_reg_reg_11_ ( .D(n857), .CK(clk), .RN(rstx), 
        .Q(ic_socket_gcu_o1_data0_wire[11]) );
  DFFRX2 fu_LSU_addr_reg_reg_12_ ( .D(n1083), .CK(clk), .RN(rstx), .Q(
        fu_LSU_addr[12]) );
  DFFRX1 fu_ALU_t1reg_reg_14_ ( .D(n1081), .CK(clk), .RN(rstx), .Q(
        fu_ALU_t1reg[14]) );
  DFFRX1 fu_ALU_t1reg_reg_16_ ( .D(n792), .CK(clk), .RN(rstx), .Q(
        fu_ALU_t1reg[16]) );
  DFFRX2 fu_LSU_data_out_reg_reg_2_ ( .D(n979), .CK(clk), .RN(rstx), .Q(
        fu_LSU_data_out[2]) );
  DFFRX2 fu_LSU_data_out_reg_reg_7_ ( .D(n904), .CK(clk), .RN(rstx), .Q(
        fu_LSU_data_out[7]) );
  DFFRX2 fu_LSU_data_out_reg_reg_6_ ( .D(n919), .CK(clk), .RN(rstx), .Q(
        fu_LSU_data_out[6]) );
  DFFRX2 fu_LSU_data_out_reg_reg_5_ ( .D(n934), .CK(clk), .RN(rstx), .Q(
        fu_LSU_data_out[5]) );
  DFFRX2 fu_LSU_data_out_reg_reg_4_ ( .D(n949), .CK(clk), .RN(rstx), .Q(
        fu_LSU_data_out[4]) );
  DFFRX2 fu_LSU_data_out_reg_reg_3_ ( .D(n964), .CK(clk), .RN(rstx), .Q(
        fu_LSU_data_out[3]) );
  DFFRX2 fu_ALU_o1temp_reg_13_ ( .D(n821), .CK(clk), .RN(rstx), .QN(n268) );
  DFFRX2 rf_RF_reg_reg_4__13_ ( .D(n826), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_4__13_) );
  DFFRX2 rf_RF_reg_reg_3__13_ ( .D(n825), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_3__13_) );
  DFFRX2 rf_RF_reg_reg_2__13_ ( .D(n824), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_2__13_) );
  DFFRX2 rf_RF_reg_reg_1__13_ ( .D(n823), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_1__13_) );
  DFFRX2 rf_RF_reg_reg_0__13_ ( .D(n822), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_0__13_) );
  DFFRX2 fu_LSU_o1shadow_reg_reg_13_ ( .D(n819), .CK(clk), .RN(rstx), .Q(
        fu_LSU_o1shadow_reg_13_) );
  DFFRX2 fu_ALU_o1temp_reg_15_ ( .D(n804), .CK(clk), .RN(rstx), .QN(n248) );
  DFFRX2 rf_RF_reg_reg_4__15_ ( .D(n809), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_4__15_) );
  DFFRX2 rf_RF_reg_reg_3__15_ ( .D(n808), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_3__15_) );
  DFFRX2 rf_RF_reg_reg_2__15_ ( .D(n807), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_2__15_) );
  DFFRX2 rf_RF_reg_reg_1__15_ ( .D(n806), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_1__15_) );
  DFFRX2 rf_RF_reg_reg_0__15_ ( .D(n805), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_0__15_) );
  DFFRX2 fu_LSU_data_out_reg_reg_13_ ( .D(n814), .CK(clk), .RN(rstx), .Q(
        fu_LSU_data_out[13]) );
  DFFRX2 fu_LSU_data_out_reg_reg_15_ ( .D(n801), .CK(clk), .RN(rstx), .Q(
        fu_LSU_data_out[15]) );
  DFFRX2 inst_fetch_return_addr_reg_reg_13_ ( .D(n827), .CK(clk), .RN(rstx), 
        .Q(ic_socket_gcu_o1_data0_wire[13]) );
  DFFRX1 fu_ALU_t1reg_reg_17_ ( .D(n782), .CK(clk), .RN(rstx), .Q(
        fu_ALU_t1reg[17]) );
  DFFRX2 rf_RF_reg_reg_4__16_ ( .D(n799), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_4__16_) );
  DFFRX2 rf_RF_reg_reg_3__16_ ( .D(n798), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_3__16_) );
  DFFRX2 rf_RF_reg_reg_2__16_ ( .D(n797), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_2__16_) );
  DFFRX2 rf_RF_reg_reg_1__16_ ( .D(n796), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_1__16_) );
  DFFRX2 rf_RF_reg_reg_0__16_ ( .D(n795), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_0__16_) );
  DFFRX2 fu_ALU_o1temp_reg_16_ ( .D(n794), .CK(clk), .RN(rstx), .QN(n228) );
  DFFRX2 fu_LSU_o1shadow_reg_reg_16_ ( .D(n793), .CK(clk), .RN(rstx), .Q(
        fu_LSU_o1shadow_reg_16_) );
  DFFRX2 rf_RF_reg_reg_4__14_ ( .D(n1089), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_4__14_) );
  DFFRX2 rf_RF_reg_reg_3__14_ ( .D(n1088), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_3__14_) );
  DFFRX2 rf_RF_reg_reg_2__14_ ( .D(n1087), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_2__14_) );
  DFFRX2 rf_RF_reg_reg_1__14_ ( .D(n1086), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_1__14_) );
  DFFRX2 rf_RF_reg_reg_0__14_ ( .D(n1085), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_0__14_) );
  DFFRX2 fu_ALU_o1temp_reg_14_ ( .D(n1084), .CK(clk), .RN(rstx), .QN(n260) );
  DFFRX2 fu_LSU_o1shadow_reg_reg_14_ ( .D(n1082), .CK(clk), .RN(rstx), .Q(
        fu_LSU_o1shadow_reg_14_) );
  DFFRX2 fu_LSU_data_out_reg_reg_14_ ( .D(n811), .CK(clk), .RN(rstx), .Q(
        fu_LSU_data_out[14]) );
  DFFRX2 inst_fetch_return_addr_reg_reg_14_ ( .D(n812), .CK(clk), .RN(rstx), 
        .Q(ic_socket_gcu_o1_data0_wire[14]) );
  DFFRX1 fu_ALU_t1reg_reg_18_ ( .D(n772), .CK(clk), .RN(rstx), .Q(
        fu_ALU_t1reg[18]) );
  DFFRX2 fu_LSU_data_out_reg_reg_17_ ( .D(n781), .CK(clk), .RN(rstx), .Q(
        fu_LSU_data_out[17]) );
  DFFRX2 rf_RF_reg_reg_4__17_ ( .D(n789), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_4__17_) );
  DFFRX2 rf_RF_reg_reg_3__17_ ( .D(n788), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_3__17_) );
  DFFRX2 rf_RF_reg_reg_2__17_ ( .D(n787), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_2__17_) );
  DFFRX2 rf_RF_reg_reg_1__17_ ( .D(n786), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_1__17_) );
  DFFRX2 rf_RF_reg_reg_0__17_ ( .D(n785), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_0__17_) );
  DFFRX2 fu_ALU_o1temp_reg_17_ ( .D(n784), .CK(clk), .RN(rstx), .QN(n215) );
  DFFRX2 fu_LSU_o1shadow_reg_reg_17_ ( .D(n783), .CK(clk), .RN(rstx), .Q(
        fu_LSU_o1shadow_reg_17_) );
  DFFRX2 fu_LSU_data_out_reg_reg_18_ ( .D(n771), .CK(clk), .RN(rstx), .Q(
        fu_LSU_data_out[18]) );
  DFFRX1 fu_ALU_t1reg_reg_19_ ( .D(n762), .CK(clk), .RN(rstx), .Q(
        fu_ALU_t1reg[19]) );
  DFFRX2 fu_LSU_data_out_reg_reg_16_ ( .D(n791), .CK(clk), .RN(rstx), .Q(
        fu_LSU_data_out[16]) );
  DFFRX2 rf_RF_reg_reg_4__18_ ( .D(n779), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_4__18_) );
  DFFRX2 rf_RF_reg_reg_3__18_ ( .D(n778), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_3__18_) );
  DFFRX2 rf_RF_reg_reg_2__18_ ( .D(n777), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_2__18_) );
  DFFRX2 rf_RF_reg_reg_1__18_ ( .D(n776), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_1__18_) );
  DFFRX2 rf_RF_reg_reg_0__18_ ( .D(n775), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_0__18_) );
  DFFRX2 fu_ALU_o1temp_reg_18_ ( .D(n774), .CK(clk), .RN(rstx), .QN(n201) );
  DFFRX2 fu_LSU_o1shadow_reg_reg_18_ ( .D(n773), .CK(clk), .RN(rstx), .Q(
        fu_LSU_o1shadow_reg_18_) );
  DFFRX2 fu_LSU_data_out_reg_reg_19_ ( .D(n761), .CK(clk), .RN(rstx), .Q(
        fu_LSU_data_out[19]) );
  DFFRX1 fu_ALU_t1reg_reg_20_ ( .D(n752), .CK(clk), .RN(rstx), .Q(
        fu_ALU_t1reg[20]) );
  DFFRX2 rf_RF_reg_reg_4__19_ ( .D(n769), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_4__19_) );
  DFFRX2 rf_RF_reg_reg_3__19_ ( .D(n768), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_3__19_) );
  DFFRX2 rf_RF_reg_reg_2__19_ ( .D(n767), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_2__19_) );
  DFFRX2 rf_RF_reg_reg_1__19_ ( .D(n766), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_1__19_) );
  DFFRX2 rf_RF_reg_reg_0__19_ ( .D(n765), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_0__19_) );
  DFFRX2 fu_ALU_o1temp_reg_19_ ( .D(n764), .CK(clk), .RN(rstx), .QN(n189) );
  DFFRX2 fu_LSU_o1shadow_reg_reg_19_ ( .D(n763), .CK(clk), .RN(rstx), .Q(
        fu_LSU_o1shadow_reg_19_) );
  DFFRX2 inst_decoder_fu_LIFTING_x2_load_reg_reg ( .D(n1145), .CK(clk), .RN(
        rstx), .Q(fu_LIFTING_in2_load_wire) );
  DFFRX2 fu_LSU_data_out_reg_reg_20_ ( .D(n751), .CK(clk), .RN(rstx), .Q(
        fu_LSU_data_out[20]) );
  DFFRX2 inst_decoder_socket_bool_o1_bus_cntrl_reg_reg_0_ ( .D(n1186), .CK(clk), .RN(rstx), .Q(ic_socket_bool_o1_bus_cntrl_wire_0_) );
  DFFRX2 fu_ALU_o1temp_reg_20_ ( .D(n754), .CK(clk), .RN(rstx), .QN(n177) );
  DFFRX2 fu_LSU_o1shadow_reg_reg_20_ ( .D(n753), .CK(clk), .RN(rstx), .Q(
        fu_LSU_o1shadow_reg_20_) );
  DFFRX2 rf_RF_reg_reg_4__20_ ( .D(n759), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_4__20_) );
  DFFRX2 rf_RF_reg_reg_3__20_ ( .D(n758), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_3__20_) );
  DFFRX2 rf_RF_reg_reg_2__20_ ( .D(n757), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_2__20_) );
  DFFRX2 rf_RF_reg_reg_1__20_ ( .D(n756), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_1__20_) );
  DFFRX2 rf_RF_reg_reg_0__20_ ( .D(n755), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_0__20_) );
  DFFRX2 fu_LSU_data_out_reg_reg_21_ ( .D(n741), .CK(clk), .RN(rstx), .Q(
        fu_LSU_data_out[21]) );
  DFFRX1 fu_ALU_t1reg_reg_22_ ( .D(n732), .CK(clk), .RN(rstx), .Q(
        fu_ALU_t1reg[22]) );
  DFFRX2 fu_ALU_o1temp_reg_21_ ( .D(n744), .CK(clk), .RN(rstx), .QN(n165) );
  DFFRX2 rf_RF_reg_reg_4__21_ ( .D(n749), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_4__21_) );
  DFFRX2 rf_RF_reg_reg_3__21_ ( .D(n748), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_3__21_) );
  DFFRX2 rf_RF_reg_reg_2__21_ ( .D(n747), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_2__21_) );
  DFFRX2 rf_RF_reg_reg_1__21_ ( .D(n746), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_1__21_) );
  DFFRX2 rf_RF_reg_reg_0__21_ ( .D(n745), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_0__21_) );
  DFFRX2 fu_LSU_o1shadow_reg_reg_21_ ( .D(n743), .CK(clk), .RN(rstx), .Q(
        fu_LSU_o1shadow_reg_21_) );
  DFFRX2 inst_decoder_simm_B1_reg_reg_26_ ( .D(n1149), .CK(clk), .RN(rstx), 
        .Q(ic_simm_B1_wire[26]) );
  DFFRX2 fu_LSU_data_out_reg_reg_22_ ( .D(n731), .CK(clk), .RN(rstx), .Q(
        fu_LSU_data_out[22]) );
  DFFRX2 inst_decoder_rf_BOOL_wr_load_reg_reg ( .D(n1138), .CK(clk), .RN(rstx), 
        .Q(rf_BOOL_t1load_wire), .QN(n561) );
  DFFRX2 rf_RF_reg_reg_4__22_ ( .D(n739), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_4__22_) );
  DFFRX2 rf_RF_reg_reg_3__22_ ( .D(n738), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_3__22_) );
  DFFRX2 rf_RF_reg_reg_2__22_ ( .D(n737), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_2__22_) );
  DFFRX2 rf_RF_reg_reg_1__22_ ( .D(n736), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_1__22_) );
  DFFRX2 rf_RF_reg_reg_0__22_ ( .D(n735), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_0__22_) );
  DFFRX2 fu_ALU_o1temp_reg_22_ ( .D(n734), .CK(clk), .RN(rstx), .QN(n153) );
  DFFRX2 fu_LSU_o1shadow_reg_reg_22_ ( .D(n733), .CK(clk), .RN(rstx), .Q(
        fu_LSU_o1shadow_reg_22_) );
  DFFRX2 inst_decoder_rf_RF_rd_opc_reg_reg_2_ ( .D(n1182), .CK(clk), .RN(rstx), 
        .Q(rf_RF_r1opcode_wire[2]), .QN(n585) );
  DFFRX2 fu_LSU_data_out_reg_reg_23_ ( .D(n721), .CK(clk), .RN(rstx), .Q(
        fu_LSU_data_out[23]) );
  DFFRX2 inst_decoder_socket_LIFTING_o1_bus_cntrl_reg_reg_0_ ( .D(n1189), .CK(
        clk), .RN(rstx), .Q(ic_socket_LIFTING_o1_bus_cntrl_wire_0_) );
  DFFRX2 inst_decoder_socket_ALU_o1_bus_cntrl_reg_reg_0_ ( .D(n1187), .CK(clk), 
        .RN(rstx), .Q(ic_socket_ALU_o1_bus_cntrl_wire_0_) );
  DFFRX2 inst_decoder_fu_ALU_in1t_load_reg_reg ( .D(n1122), .CK(clk), .RN(rstx), .Q(fu_ALU_t1load_wire) );
  DFFRX2 inst_decoder_fu_gcu_opc_reg_reg_0_ ( .D(n1134), .CK(clk), .RN(rstx), 
        .Q(inst_fetch_pc_opcode_wire_0_) );
  DFFRX1 fu_ALU_t1reg_reg_24_ ( .D(n712), .CK(clk), .RN(rstx), .Q(
        fu_ALU_t1reg[24]) );
  DFFRX2 fu_ALU_o1temp_reg_23_ ( .D(n724), .CK(clk), .RN(rstx), .QN(n139) );
  DFFRX2 fu_LSU_o1shadow_reg_reg_23_ ( .D(n723), .CK(clk), .RN(rstx), .Q(
        fu_LSU_o1shadow_reg_23_) );
  DFFRX2 rf_RF_reg_reg_4__23_ ( .D(n729), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_4__23_) );
  DFFRX2 rf_RF_reg_reg_3__23_ ( .D(n728), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_3__23_) );
  DFFRX2 rf_RF_reg_reg_2__23_ ( .D(n727), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_2__23_) );
  DFFRX2 rf_RF_reg_reg_1__23_ ( .D(n726), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_1__23_) );
  DFFRX2 rf_RF_reg_reg_0__23_ ( .D(n725), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_0__23_) );
  DFFRX1 inst_decoder_socket_gcu_o1_bus_cntrl_reg_reg_0_ ( .D(n1184), .CK(clk), 
        .RN(rstx), .Q(ic_socket_gcu_o1_bus_cntrl_wire_0_) );
  DFFRX2 inst_decoder_simm_B1_reg_reg_1_ ( .D(n1163), .CK(clk), .RN(rstx), .Q(
        ic_simm_B1_wire[1]) );
  DFFRX2 inst_decoder_fu_ALU_opc_reg_reg_3_ ( .D(n1120), .CK(clk), .RN(rstx), 
        .Q(fu_ALU_t1opcode_wire[3]) );
  DFFRX2 inst_decoder_fu_ALU_opc_reg_reg_0_ ( .D(n1116), .CK(clk), .RN(rstx), 
        .Q(fu_ALU_t1opcode_wire[0]) );
  DFFRX2 inst_decoder_fu_ALU_opc_reg_reg_1_ ( .D(n1118), .CK(clk), .RN(rstx), 
        .Q(fu_ALU_t1opcode_wire[1]) );
  DFFRX2 inst_decoder_fu_ALU_opc_reg_reg_2_ ( .D(n1114), .CK(clk), .RN(rstx), 
        .Q(fu_ALU_t1opcode_wire[2]) );
  DFFRX2 inst_decoder_simm_B1_reg_reg_2_ ( .D(n1161), .CK(clk), .RN(rstx), .Q(
        ic_simm_B1_wire[2]) );
  DFFRX2 inst_decoder_simm_B1_reg_reg_0_ ( .D(n1162), .CK(clk), .RN(rstx), .Q(
        ic_simm_B1_wire[0]) );
  DFFRX2 inst_decoder_rf_RF_wr_load_reg_reg ( .D(n1131), .CK(clk), .RN(rstx), 
        .Q(rf_RF_t1load_wire) );
  DFFRX2 fu_LSU_data_out_reg_reg_24_ ( .D(n711), .CK(clk), .RN(rstx), .Q(
        fu_LSU_data_out[24]) );
  DFFRX1 fu_ALU_t1reg_reg_25_ ( .D(n702), .CK(clk), .RN(rstx), .Q(
        fu_ALU_t1reg[25]) );
  DFFRX2 rf_RF_reg_reg_4__24_ ( .D(n719), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_4__24_) );
  DFFRX2 rf_RF_reg_reg_3__24_ ( .D(n718), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_3__24_) );
  DFFRX2 rf_RF_reg_reg_2__24_ ( .D(n717), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_2__24_) );
  DFFRX2 rf_RF_reg_reg_1__24_ ( .D(n716), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_1__24_) );
  DFFRX2 rf_RF_reg_reg_0__24_ ( .D(n715), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_0__24_) );
  DFFRX2 fu_ALU_o1temp_reg_24_ ( .D(n714), .CK(clk), .RN(rstx), .QN(n123) );
  DFFRX2 fu_LSU_o1shadow_reg_reg_24_ ( .D(n713), .CK(clk), .RN(rstx), .Q(
        fu_LSU_o1shadow_reg_24_) );
  DFFRX1 fu_ALU_t1reg_reg_26_ ( .D(n692), .CK(clk), .RN(rstx), .Q(
        fu_ALU_t1reg[26]) );
  DFFRX2 rf_RF_reg_reg_4__25_ ( .D(n709), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_4__25_) );
  DFFRX2 rf_RF_reg_reg_3__25_ ( .D(n708), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_3__25_) );
  DFFRX2 rf_RF_reg_reg_2__25_ ( .D(n707), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_2__25_) );
  DFFRX2 rf_RF_reg_reg_1__25_ ( .D(n706), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_1__25_) );
  DFFRX2 rf_RF_reg_reg_0__25_ ( .D(n705), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_0__25_) );
  DFFRX2 fu_ALU_o1temp_reg_25_ ( .D(n704), .CK(clk), .RN(rstx), .QN(n110) );
  DFFRX2 fu_LSU_o1shadow_reg_reg_25_ ( .D(n703), .CK(clk), .RN(rstx), .Q(
        fu_LSU_o1shadow_reg_25_) );
  DFFRX2 inst_decoder_simm_B1_reg_reg_28_ ( .D(n1148), .CK(clk), .RN(rstx), 
        .Q(ic_simm_B1_wire[28]) );
  DFFRX2 inst_decoder_simm_B1_reg_reg_27_ ( .D(n1176), .CK(clk), .RN(rstx), 
        .Q(ic_simm_B1_wire[27]) );
  DFFRX2 inst_decoder_simm_B1_reg_reg_25_ ( .D(n1175), .CK(clk), .RN(rstx), 
        .Q(ic_simm_B1_wire[25]) );
  DFFRX2 inst_decoder_simm_B1_reg_reg_24_ ( .D(n1150), .CK(clk), .RN(rstx), 
        .Q(ic_simm_B1_wire[24]) );
  DFFRX2 inst_decoder_simm_B1_reg_reg_23_ ( .D(n1174), .CK(clk), .RN(rstx), 
        .Q(ic_simm_B1_wire[23]) );
  DFFRX2 inst_decoder_simm_B1_reg_reg_22_ ( .D(n1151), .CK(clk), .RN(rstx), 
        .Q(ic_simm_B1_wire[22]) );
  DFFRX2 inst_decoder_simm_B1_reg_reg_21_ ( .D(n1173), .CK(clk), .RN(rstx), 
        .Q(ic_simm_B1_wire[21]) );
  DFFRX2 inst_decoder_simm_B1_reg_reg_20_ ( .D(n1152), .CK(clk), .RN(rstx), 
        .Q(ic_simm_B1_wire[20]) );
  DFFRX2 inst_decoder_simm_B1_reg_reg_19_ ( .D(n1172), .CK(clk), .RN(rstx), 
        .Q(ic_simm_B1_wire[19]) );
  DFFRX2 inst_decoder_simm_B1_reg_reg_18_ ( .D(n1153), .CK(clk), .RN(rstx), 
        .Q(ic_simm_B1_wire[18]) );
  DFFRX2 inst_decoder_simm_B1_reg_reg_17_ ( .D(n1171), .CK(clk), .RN(rstx), 
        .Q(ic_simm_B1_wire[17]) );
  DFFRX2 inst_decoder_simm_B1_reg_reg_16_ ( .D(n1154), .CK(clk), .RN(rstx), 
        .Q(ic_simm_B1_wire[16]) );
  DFFRX2 inst_decoder_simm_B1_reg_reg_15_ ( .D(n1170), .CK(clk), .RN(rstx), 
        .Q(ic_simm_B1_wire[15]) );
  DFFRX2 inst_decoder_simm_B1_reg_reg_14_ ( .D(n1155), .CK(clk), .RN(rstx), 
        .Q(ic_simm_B1_wire[14]) );
  DFFRX2 inst_decoder_simm_B1_reg_reg_13_ ( .D(n1169), .CK(clk), .RN(rstx), 
        .Q(ic_simm_B1_wire[13]) );
  DFFRX2 inst_decoder_simm_B1_reg_reg_12_ ( .D(n1156), .CK(clk), .RN(rstx), 
        .Q(ic_simm_B1_wire[12]) );
  DFFRX2 inst_decoder_simm_B1_reg_reg_11_ ( .D(n1168), .CK(clk), .RN(rstx), 
        .Q(ic_simm_B1_wire[11]) );
  DFFRX2 inst_decoder_simm_B1_reg_reg_10_ ( .D(n1157), .CK(clk), .RN(rstx), 
        .Q(ic_simm_B1_wire[10]) );
  DFFRX2 inst_decoder_simm_B1_reg_reg_9_ ( .D(n1167), .CK(clk), .RN(rstx), .Q(
        ic_simm_B1_wire[9]) );
  DFFRX2 inst_decoder_simm_B1_reg_reg_8_ ( .D(n1158), .CK(clk), .RN(rstx), .Q(
        ic_simm_B1_wire[8]) );
  DFFRX2 inst_decoder_simm_B1_reg_reg_7_ ( .D(n1166), .CK(clk), .RN(rstx), .Q(
        ic_simm_B1_wire[7]) );
  DFFRX2 inst_decoder_simm_B1_reg_reg_6_ ( .D(n1159), .CK(clk), .RN(rstx), .Q(
        ic_simm_B1_wire[6]) );
  DFFRX2 inst_decoder_simm_B1_reg_reg_5_ ( .D(n1165), .CK(clk), .RN(rstx), .Q(
        ic_simm_B1_wire[5]) );
  DFFRX2 inst_decoder_simm_B1_reg_reg_4_ ( .D(n1160), .CK(clk), .RN(rstx), .Q(
        ic_simm_B1_wire[4]) );
  DFFRX2 inst_decoder_simm_B1_reg_reg_3_ ( .D(n1164), .CK(clk), .RN(rstx), .Q(
        ic_simm_B1_wire[3]) );
  DFFRX2 inst_decoder_simm_B1_reg_reg_30_ ( .D(n1147), .CK(clk), .RN(rstx), 
        .QN(n49) );
  DFFRX2 inst_decoder_simm_B1_reg_reg_31_ ( .D(n1178), .CK(clk), .RN(rstx), 
        .QN(n513) );
  DFFRX2 inst_decoder_simm_B1_reg_reg_29_ ( .D(n1177), .CK(clk), .RN(rstx), 
        .QN(n67) );
  DFFRX2 fu_LSU_data_out_reg_reg_25_ ( .D(n701), .CK(clk), .RN(rstx), .Q(
        fu_LSU_data_out[25]) );
  DFFRX2 fu_LSU_data_out_reg_reg_26_ ( .D(n691), .CK(clk), .RN(rstx), .Q(
        fu_LSU_data_out[26]) );
  DFFRX1 fu_ALU_t1reg_reg_27_ ( .D(n682), .CK(clk), .RN(rstx), .Q(
        fu_ALU_t1reg[27]) );
  DFFRX2 rf_RF_reg_reg_4__26_ ( .D(n699), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_4__26_) );
  DFFRX2 rf_RF_reg_reg_3__26_ ( .D(n698), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_3__26_) );
  DFFRX2 rf_RF_reg_reg_2__26_ ( .D(n697), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_2__26_) );
  DFFRX2 rf_RF_reg_reg_1__26_ ( .D(n696), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_1__26_) );
  DFFRX2 rf_RF_reg_reg_0__26_ ( .D(n695), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_0__26_) );
  DFFRX2 fu_ALU_o1temp_reg_26_ ( .D(n694), .CK(clk), .RN(rstx), .QN(n97) );
  DFFRX2 fu_LSU_o1shadow_reg_reg_26_ ( .D(n693), .CK(clk), .RN(rstx), .Q(
        fu_LSU_o1shadow_reg_26_) );
  DFFRX2 fu_LSU_data_out_reg_reg_27_ ( .D(n681), .CK(clk), .RN(rstx), .Q(
        fu_LSU_data_out[27]) );
  DFFRX2 rf_RF_reg_reg_4__27_ ( .D(n689), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_4__27_) );
  DFFRX2 rf_RF_reg_reg_3__27_ ( .D(n688), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_3__27_) );
  DFFRX2 rf_RF_reg_reg_2__27_ ( .D(n687), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_2__27_) );
  DFFRX2 rf_RF_reg_reg_1__27_ ( .D(n686), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_1__27_) );
  DFFRX2 rf_RF_reg_reg_0__27_ ( .D(n685), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_0__27_) );
  DFFRX2 fu_ALU_o1temp_reg_27_ ( .D(n684), .CK(clk), .RN(rstx), .QN(n85) );
  DFFRX2 fu_LSU_o1shadow_reg_reg_27_ ( .D(n683), .CK(clk), .RN(rstx), .Q(
        fu_LSU_o1shadow_reg_27_) );
  DFFRX1 fu_ALU_o1reg_reg_27_ ( .D(n680), .CK(clk), .RN(rstx), .Q(
        fu_ALU_o1reg[27]) );
  DFFRX2 fu_LSU_data_out_reg_reg_28_ ( .D(n671), .CK(clk), .RN(rstx), .Q(
        fu_LSU_data_out[28]) );
  DFFRX1 fu_ALU_t1reg_reg_29_ ( .D(n662), .CK(clk), .RN(rstx), .Q(
        fu_ALU_t1reg[29]) );
  DFFRX2 rf_RF_reg_reg_4__28_ ( .D(n679), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_4__28_) );
  DFFRX2 rf_RF_reg_reg_3__28_ ( .D(n678), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_3__28_) );
  DFFRX2 rf_RF_reg_reg_2__28_ ( .D(n677), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_2__28_) );
  DFFRX2 rf_RF_reg_reg_1__28_ ( .D(n676), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_1__28_) );
  DFFRX2 rf_RF_reg_reg_0__28_ ( .D(n675), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_0__28_) );
  DFFRX2 fu_ALU_o1temp_reg_28_ ( .D(n674), .CK(clk), .RN(rstx), .QN(n73) );
  DFFRX2 fu_LSU_o1shadow_reg_reg_28_ ( .D(n673), .CK(clk), .RN(rstx), .Q(
        fu_LSU_o1shadow_reg_28_) );
  DFFRX2 fu_LSU_data_out_reg_reg_29_ ( .D(n661), .CK(clk), .RN(rstx), .Q(
        fu_LSU_data_out[29]) );
  DFFRX2 rf_RF_reg_reg_4__29_ ( .D(n669), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_4__29_) );
  DFFRX2 rf_RF_reg_reg_3__29_ ( .D(n668), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_3__29_) );
  DFFRX2 rf_RF_reg_reg_2__29_ ( .D(n667), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_2__29_) );
  DFFRX2 rf_RF_reg_reg_1__29_ ( .D(n666), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_1__29_) );
  DFFRX2 rf_RF_reg_reg_0__29_ ( .D(n665), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_0__29_) );
  DFFRX2 fu_ALU_o1temp_reg_29_ ( .D(n664), .CK(clk), .RN(rstx), .QN(n60) );
  DFFRX2 fu_LSU_o1shadow_reg_reg_29_ ( .D(n663), .CK(clk), .RN(rstx), .Q(
        fu_LSU_o1shadow_reg_29_) );
  DFFRX1 fu_ALU_t1reg_reg_30_ ( .D(n652), .CK(clk), .RN(rstx), .Q(
        fu_ALU_t1reg[30]) );
  DFFRX2 fu_LSU_data_out_reg_reg_30_ ( .D(n651), .CK(clk), .RN(rstx), .Q(
        fu_LSU_data_out[30]) );
  DFFRX2 fu_LSU_data_out_reg_reg_31_ ( .D(n649), .CK(clk), .RN(rstx), .Q(
        fu_LSU_data_out[31]) );
  DFFRX2 rf_RF_reg_reg_4__30_ ( .D(n659), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_4__30_) );
  DFFRX2 rf_RF_reg_reg_3__30_ ( .D(n658), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_3__30_) );
  DFFRX2 rf_RF_reg_reg_2__30_ ( .D(n657), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_2__30_) );
  DFFRX2 rf_RF_reg_reg_1__30_ ( .D(n656), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_1__30_) );
  DFFRX2 rf_RF_reg_reg_0__30_ ( .D(n655), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_0__30_) );
  DFFRX2 fu_ALU_o1temp_reg_30_ ( .D(n654), .CK(clk), .RN(rstx), .QN(n33) );
  DFFRX2 fu_LSU_o1shadow_reg_reg_30_ ( .D(n653), .CK(clk), .RN(rstx), .Q(
        fu_LSU_o1shadow_reg_30_) );
  DFFRX2 rf_RF_reg_reg_4__31_ ( .D(n1097), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_4__31_) );
  DFFRX2 rf_RF_reg_reg_3__31_ ( .D(n1096), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_3__31_) );
  DFFRX2 rf_RF_reg_reg_2__31_ ( .D(n1095), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_2__31_) );
  DFFRX2 rf_RF_reg_reg_1__31_ ( .D(n1094), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_1__31_) );
  DFFRX2 rf_RF_reg_reg_0__31_ ( .D(n1093), .CK(clk), .RN(rstx), .Q(
        rf_RF_reg_0__31_) );
  DFFRX2 fu_ALU_o1temp_reg_31_ ( .D(n1092), .CK(clk), .RN(rstx), .QN(n20) );
  DFFRX2 fu_LSU_o1shadow_reg_reg_31_ ( .D(n1091), .CK(clk), .RN(rstx), .Q(
        fu_LSU_o1shadow_reg_31_) );
  OR2X2 U1284 ( .A(n2249), .B(n1286), .Y(n1267) );
  INVX5 U1285 ( .A(n1267), .Y(n1268) );
  OR3X2 U1286 ( .A(n2183), .B(n2111), .C(n2249), .Y(n1269) );
  CLKINVX4 U1287 ( .A(n1269), .Y(n1270) );
  OR2XL U1288 ( .A(n1268), .B(n1826), .Y(n1271) );
  CLKINVX8 U1289 ( .A(n1271), .Y(n1272) );
  OR2XL U1290 ( .A(n1270), .B(n1826), .Y(n1273) );
  CLKINVX8 U1291 ( .A(n1273), .Y(n1274) );
  OR2XL U1292 ( .A(n1270), .B(n1782), .Y(n1275) );
  CLKINVX8 U1293 ( .A(n1275), .Y(n1276) );
  OR2XL U1294 ( .A(n1268), .B(n1782), .Y(n1277) );
  CLKINVX8 U1295 ( .A(n1277), .Y(n1278) );
  OR3X2 U1296 ( .A(n452), .B(fu_LSU_status_addr_reg_1__1_), .C(n2212), .Y(
        n1279) );
  CLKINVX8 U1297 ( .A(n1279), .Y(n1280) );
  AND2X2 U1298 ( .A(inst_fetch_pc_load_wire), .B(n2208), .Y(n1281) );
  INVX14 U1299 ( .A(n1281), .Y(n1282) );
  AO22X1 U1300 ( .A0(n206), .A1(n332), .B0(n2110), .B1(n1268), .Y(n1283) );
  INVX5 U1301 ( .A(n1283), .Y(n1284) );
  BUFX12 U1302 ( .A(n2097), .Y(n1285) );
  NOR2BX1 U1303 ( .AN(n2210), .B(n521), .Y(n2097) );
  NOR2X6 U1304 ( .A(n417), .B(n418), .Y(n206) );
  MXI2X4 U1305 ( .A(n1306), .B(n1307), .S0(n2208), .Y(imem_addr[7]) );
  MXI2X4 U1306 ( .A(n1292), .B(n1293), .S0(n2209), .Y(imem_addr[8]) );
  MXI2X4 U1307 ( .A(n1304), .B(n1305), .S0(n2208), .Y(imem_addr[6]) );
  MXI2X4 U1308 ( .A(n1308), .B(n1309), .S0(n2208), .Y(imem_addr[9]) );
  MXI2X4 U1309 ( .A(n1302), .B(n1303), .S0(n2208), .Y(imem_addr[5]) );
  MXI2X4 U1310 ( .A(n1310), .B(n1311), .S0(n2208), .Y(imem_addr[10]) );
  MXI2X4 U1311 ( .A(n1300), .B(n1301), .S0(n2208), .Y(imem_addr[4]) );
  MXI2X4 U1312 ( .A(n1312), .B(n1313), .S0(n2208), .Y(imem_addr[11]) );
  MXI2X4 U1313 ( .A(n1298), .B(n1299), .S0(n2208), .Y(imem_addr[3]) );
  MXI2X4 U1314 ( .A(n1314), .B(n1315), .S0(n2208), .Y(imem_addr[12]) );
  MXI2X4 U1315 ( .A(n1296), .B(n1297), .S0(n2208), .Y(imem_addr[2]) );
  MXI2X4 U1316 ( .A(n1316), .B(n1317), .S0(n2208), .Y(imem_addr[13]) );
  MXI2X4 U1317 ( .A(n1294), .B(n1295), .S0(n2208), .Y(imem_addr[1]) );
  MXI2X4 U1318 ( .A(n1318), .B(n1319), .S0(n2208), .Y(imem_addr[14]) );
  MXI2X4 U1319 ( .A(n1291), .B(inst_fetch_increased_pc_0_), .S0(n2209), .Y(
        imem_addr[0]) );
  NOR2X6 U1320 ( .A(n1288), .B(n1289), .Y(n1893) );
  INVX5 U1321 ( .A(n250), .Y(n332) );
  OR2X8 U1322 ( .A(n1898), .B(n2118), .Y(n1287) );
  CLKBUFX20 U1323 ( .A(n1285), .Y(n1761) );
  CLKINVX40 U1324 ( .A(n2213), .Y(n2212) );
  CLKINVX16 U1325 ( .A(n1285), .Y(n2244) );
  CLKINVX16 U1326 ( .A(n1285), .Y(n2243) );
  CLKBUFX40 U1327 ( .A(n504), .Y(n2208) );
  INVX2 U1328 ( .A(n2108), .Y(fu_ALU_fu_arch_n284) );
  NAND2X2 U1329 ( .A(n1897), .B(n2111), .Y(n1286) );
  INVX4 U1330 ( .A(busy), .Y(n504) );
  NAND2X2 U1331 ( .A(n1894), .B(inst_decoder_instructionword_wire[38]), .Y(
        n1288) );
  NAND2X2 U1332 ( .A(n1895), .B(n1896), .Y(n1289) );
  AND2X2 U1333 ( .A(n1290), .B(n494), .Y(n1900) );
  OR2X2 U1334 ( .A(n454), .B(n1901), .Y(n1290) );
  BUFX8 U1335 ( .A(fu_ALU_o1reg[0]), .Y(n2181) );
  INVX8 U1336 ( .A(n2175), .Y(fu_ALU_fu_arch_sub_200_B_2_) );
  BUFX8 U1337 ( .A(fu_ALU_o1reg[9]), .Y(fu_ALU_fu_arch_sub_200_B_9_) );
  INVX12 U1338 ( .A(n2184), .Y(n1779) );
  CLKBUFX6 U1339 ( .A(fu_ALU_fu_arch_n266), .Y(n1850) );
  CLKAND2X8 U1340 ( .A(fu_ALU_opc1reg[2]), .B(fu_ALU_opc1reg[3]), .Y(
        fu_ALU_fu_arch_n175) );
  OR4X2 U1341 ( .A(n1320), .B(n1321), .C(n1322), .D(n1323), .Y(n619) );
  OR4X2 U1342 ( .A(inst_fetch_reset_cntr_24_), .B(inst_fetch_reset_cntr_23_), 
        .C(inst_fetch_reset_cntr_20_), .D(inst_fetch_reset_cntr_22_), .Y(n1320) );
  OR4X2 U1343 ( .A(inst_fetch_reset_cntr_28_), .B(inst_fetch_reset_cntr_27_), 
        .C(inst_fetch_reset_cntr_26_), .D(inst_fetch_reset_cntr_25_), .Y(n1321) );
  OR4X2 U1344 ( .A(inst_fetch_reset_cntr_17_), .B(inst_fetch_reset_cntr_16_), 
        .C(inst_fetch_reset_cntr_15_), .D(inst_fetch_reset_cntr_14_), .Y(n1322) );
  OR4X2 U1345 ( .A(inst_fetch_reset_cntr_21_), .B(inst_fetch_reset_cntr_1_), 
        .C(inst_fetch_reset_cntr_19_), .D(inst_fetch_reset_cntr_18_), .Y(n1323) );
  NAND2BX2 U1346 ( .AN(n1324), .B(n625), .Y(n618) );
  OR4X2 U1347 ( .A(busy), .B(inst_fetch_reset_cntr_7_), .C(
        inst_fetch_reset_cntr_9_), .D(inst_fetch_reset_cntr_8_), .Y(n1324) );
  CLKXOR2X2 U1348 ( .A(fu_ALU_fu_arch_sub_200_B_29_), .B(n2128), .Y(n1920) );
  ADDFX1 U1349 ( .A(n2137), .B(fu_ALU_fu_arch_sub_200_B_not_24_), .CI(
        fu_ALU_fu_arch_sub_200_carry_24_), .CO(
        fu_ALU_fu_arch_sub_200_carry_25_), .S(fu_ALU_fu_arch_N636) );
  ADDFX1 U1350 ( .A(n2139), .B(fu_ALU_fu_arch_sub_200_B_not_23_), .CI(
        fu_ALU_fu_arch_sub_200_carry_23_), .CO(
        fu_ALU_fu_arch_sub_200_carry_24_), .S(fu_ALU_fu_arch_N635) );
  ADDFX1 U1351 ( .A(n2141), .B(fu_ALU_fu_arch_sub_200_B_not_22_), .CI(
        fu_ALU_fu_arch_sub_200_carry_22_), .CO(
        fu_ALU_fu_arch_sub_200_carry_23_), .S(fu_ALU_fu_arch_N634) );
  ADDFX1 U1352 ( .A(n2141), .B(fu_ALU_o1reg[22]), .CI(
        fu_ALU_fu_arch_add_171_carry_22_), .CO(
        fu_ALU_fu_arch_add_171_carry_23_), .S(fu_ALU_fu_arch_N55) );
  ADDFX1 U1353 ( .A(n2143), .B(fu_ALU_fu_arch_sub_200_B_not_21_), .CI(
        fu_ALU_fu_arch_sub_200_carry_21_), .CO(
        fu_ALU_fu_arch_sub_200_carry_22_), .S(fu_ALU_fu_arch_N633) );
  ADDFX1 U1354 ( .A(n2145), .B(fu_ALU_fu_arch_sub_200_B_not_20_), .CI(
        fu_ALU_fu_arch_sub_200_carry_20_), .CO(
        fu_ALU_fu_arch_sub_200_carry_21_), .S(fu_ALU_fu_arch_N632) );
  ADDFX1 U1355 ( .A(n2145), .B(fu_ALU_o1reg[20]), .CI(
        fu_ALU_fu_arch_add_171_carry_20_), .CO(
        fu_ALU_fu_arch_add_171_carry_21_), .S(fu_ALU_fu_arch_N53) );
  ADDFX1 U1356 ( .A(n2147), .B(n2146), .CI(fu_ALU_fu_arch_sub_200_carry_19_), 
        .CO(fu_ALU_fu_arch_sub_200_carry_20_), .S(fu_ALU_fu_arch_N631) );
  ADDFX1 U1357 ( .A(n2147), .B(fu_ALU_fu_arch_sub_200_B_19_), .CI(
        fu_ALU_fu_arch_add_171_carry_19_), .CO(
        fu_ALU_fu_arch_add_171_carry_20_), .S(fu_ALU_fu_arch_N52) );
  ADDFX1 U1358 ( .A(n2149), .B(fu_ALU_fu_arch_sub_200_B_18_), .CI(
        fu_ALU_fu_arch_add_171_carry_18_), .CO(
        fu_ALU_fu_arch_add_171_carry_19_), .S(fu_ALU_fu_arch_N51) );
  ADDFX1 U1359 ( .A(n2149), .B(n1771), .CI(fu_ALU_fu_arch_sub_200_carry_18_), 
        .CO(fu_ALU_fu_arch_sub_200_carry_19_), .S(fu_ALU_fu_arch_N630) );
  ADDFX1 U1360 ( .A(n2150), .B(fu_ALU_fu_arch_sub_200_B_not_17_), .CI(
        fu_ALU_fu_arch_sub_200_carry_17_), .CO(
        fu_ALU_fu_arch_sub_200_carry_18_), .S(fu_ALU_fu_arch_N629) );
  ADDFX1 U1361 ( .A(n2152), .B(fu_ALU_fu_arch_sub_200_B_not_16_), .CI(
        fu_ALU_fu_arch_sub_200_carry_16_), .CO(
        fu_ALU_fu_arch_sub_200_carry_17_), .S(fu_ALU_fu_arch_N628) );
  ADDFX1 U1362 ( .A(n2154), .B(n1746), .CI(fu_ALU_fu_arch_sub_200_carry_15_), 
        .CO(fu_ALU_fu_arch_sub_200_carry_16_), .S(fu_ALU_fu_arch_N627) );
  ADDFX1 U1363 ( .A(n2135), .B(n2134), .CI(fu_ALU_fu_arch_sub_200_carry_25_), 
        .CO(fu_ALU_fu_arch_sub_200_carry_26_), .S(fu_ALU_fu_arch_N637) );
  ADDFX1 U1364 ( .A(n2150), .B(fu_ALU_o1reg[17]), .CI(
        fu_ALU_fu_arch_add_171_carry_17_), .CO(
        fu_ALU_fu_arch_add_171_carry_18_), .S(fu_ALU_fu_arch_N50) );
  ADDFX1 U1365 ( .A(n2152), .B(fu_ALU_o1reg[16]), .CI(
        fu_ALU_fu_arch_add_171_carry_16_), .CO(
        fu_ALU_fu_arch_add_171_carry_17_), .S(fu_ALU_fu_arch_N49) );
  ADDFX1 U1366 ( .A(n2154), .B(n2153), .CI(fu_ALU_fu_arch_add_171_carry_15_), 
        .CO(fu_ALU_fu_arch_add_171_carry_16_), .S(fu_ALU_fu_arch_N48) );
  ADDFX1 U1367 ( .A(n2179), .B(n2155), .CI(fu_ALU_fu_arch_sub_200_carry_14_), 
        .CO(fu_ALU_fu_arch_sub_200_carry_15_), .S(fu_ALU_fu_arch_N626) );
  ADDFX1 U1368 ( .A(n2179), .B(fu_ALU_o1reg[14]), .CI(
        fu_ALU_fu_arch_add_171_carry_14_), .CO(
        fu_ALU_fu_arch_add_171_carry_15_), .S(fu_ALU_fu_arch_N47) );
  ADDFX1 U1369 ( .A(n2156), .B(fu_ALU_fu_arch_n621), .CI(
        fu_ALU_fu_arch_sub_200_carry_13_), .CO(
        fu_ALU_fu_arch_sub_200_carry_14_), .S(fu_ALU_fu_arch_N625) );
  ADDFX1 U1370 ( .A(n2158), .B(fu_ALU_fu_arch_sub_200_B_not_12_), .CI(
        fu_ALU_fu_arch_sub_200_carry_12_), .CO(
        fu_ALU_fu_arch_sub_200_carry_13_), .S(fu_ALU_fu_arch_N624) );
  ADDFX1 U1371 ( .A(n2160), .B(fu_ALU_o1reg[11]), .CI(
        fu_ALU_fu_arch_add_171_carry_11_), .CO(
        fu_ALU_fu_arch_add_171_carry_12_), .S(fu_ALU_fu_arch_N44) );
  ADDFX1 U1372 ( .A(n2163), .B(n1778), .CI(fu_ALU_fu_arch_sub_200_carry_9_), 
        .CO(fu_ALU_fu_arch_sub_200_carry_10_), .S(fu_ALU_fu_arch_N621) );
  ADDFX1 U1373 ( .A(n2156), .B(fu_ALU_o1reg[13]), .CI(
        fu_ALU_fu_arch_add_171_carry_13_), .CO(
        fu_ALU_fu_arch_add_171_carry_14_), .S(fu_ALU_fu_arch_N46) );
  ADDFX1 U1374 ( .A(n2158), .B(fu_ALU_o1reg[12]), .CI(
        fu_ALU_fu_arch_add_171_carry_12_), .CO(
        fu_ALU_fu_arch_add_171_carry_13_), .S(fu_ALU_fu_arch_N45) );
  ADDFX1 U1375 ( .A(n2160), .B(n2159), .CI(fu_ALU_fu_arch_sub_200_carry_11_), 
        .CO(fu_ALU_fu_arch_sub_200_carry_12_), .S(fu_ALU_fu_arch_N623) );
  ADDFX1 U1376 ( .A(n2162), .B(n1772), .CI(fu_ALU_fu_arch_sub_200_carry_10_), 
        .CO(fu_ALU_fu_arch_sub_200_carry_11_), .S(fu_ALU_fu_arch_N622) );
  NAND2X2 U1377 ( .A(n1779), .B(n1770), .Y(fu_ALU_fu_arch_n281) );
  NAND2BX1 U1378 ( .AN(n2204), .B(inst_fetch_add_113_carry_31_), .Y(n1734) );
  XNOR2X1 U1379 ( .A(n1734), .B(inst_fetch_reset_cntr_31_), .Y(n1265) );
  NAND2BX1 U1380 ( .AN(rstx), .B(pc_init[13]), .Y(n816) );
  NAND2BX1 U1381 ( .AN(rstx), .B(pc_init[11]), .Y(n846) );
  NAND2BX1 U1382 ( .AN(rstx), .B(pc_init[12]), .Y(n831) );
  NAND2BX1 U1383 ( .AN(rstx), .B(pc_init[10]), .Y(n861) );
  NAND2BX1 U1384 ( .AN(rstx), .B(pc_init[9]), .Y(n876) );
  NAND2BX1 U1385 ( .AN(rstx), .B(pc_init[8]), .Y(n891) );
  NAND2BX1 U1386 ( .AN(rstx), .B(pc_init[7]), .Y(n906) );
  NAND2BX1 U1387 ( .AN(rstx), .B(pc_init[6]), .Y(n921) );
  XNOR2X1 U1388 ( .A(inst_fetch_reset_cntr_0_), .B(n2205), .Y(n1248) );
  NAND4X1 U1389 ( .A(n579), .B(inst_decoder_instructionword_wire[36]), .C(
        inst_decoder_instructionword_wire[35]), .D(
        inst_decoder_instructionword_wire[38]), .Y(n1735) );
  OAI22X1 U1390 ( .A0(n1856), .A1(n1735), .B0(n149), .B1(n498), .Y(n1188) );
  OAI211X4 U1391 ( .A0(fu_ALU_fu_arch_n741), .A1(n1797), .B0(
        fu_ALU_fu_arch_n742), .C0(fu_ALU_fu_arch_n743), .Y(fu_ALU_fu_arch_n740) );
  CLKBUFX40 U1392 ( .A(rf_RF_t1data_wire[0]), .Y(n2111) );
  BUFX8 U1393 ( .A(fu_ALU_t1reg[21]), .Y(n2143) );
  BUFX8 U1394 ( .A(fu_ALU_t1reg[23]), .Y(n2139) );
  BUFX10 U1395 ( .A(fu_ALU_o1reg[1]), .Y(n2177) );
  BUFX8 U1396 ( .A(fu_ALU_t1reg[31]), .Y(n2180) );
  BUFX8 U1397 ( .A(fu_ALU_t1reg[13]), .Y(n2156) );
  INVX8 U1398 ( .A(n1753), .Y(n1754) );
  CLKBUFX16 U1399 ( .A(fu_ALU_fu_arch_n250), .Y(n2199) );
  BUFX8 U1400 ( .A(fu_ALU_t1reg[6]), .Y(n2169) );
  BUFX8 U1401 ( .A(fu_ALU_t1reg[8]), .Y(n2165) );
  BUFX8 U1402 ( .A(fu_ALU_t1reg[12]), .Y(n2158) );
  BUFX8 U1403 ( .A(fu_ALU_t1reg[9]), .Y(n2163) );
  INVX8 U1404 ( .A(n2159), .Y(fu_ALU_fu_arch_sub_200_B_11_) );
  INVX10 U1405 ( .A(n2155), .Y(fu_ALU_fu_arch_sub_200_B_14_) );
  CLKINVX8 U1406 ( .A(n2134), .Y(n1780) );
  BUFX8 U1407 ( .A(fu_ALU_t1reg[28]), .Y(n2130) );
  INVX2 U1408 ( .A(inst_decoder_instructionword_wire[38]), .Y(n580) );
  CLKXOR2X2 U1409 ( .A(n2181), .B(n1779), .Y(fu_ALU_fu_arch_N33) );
  CLKXOR2X2 U1410 ( .A(fu_ALU_fu_arch_sub_200_B_11_), .B(n2160), .Y(n1923) );
  CLKXOR2X2 U1411 ( .A(n1780), .B(n2135), .Y(n1913) );
  CLKXOR2X2 U1412 ( .A(fu_ALU_fu_arch_sub_200_B_4_), .B(n2172), .Y(n1909) );
  INVX4 U1413 ( .A(ic_socket_RF_o1_bus_cntrl_wire_0_), .Y(n1748) );
  CLKINVX3 U1414 ( .A(n1779), .Y(n1749) );
  INVX4 U1415 ( .A(ic_simm_cntrl_B1_wire_0_), .Y(n1750) );
  CLKINVX2 U1416 ( .A(n2183), .Y(n1751) );
  INVX16 U1417 ( .A(n2182), .Y(n2183) );
  INVX2 U1418 ( .A(inst_decoder_N119), .Y(n1752) );
  CLKINVX2 U1419 ( .A(n2170), .Y(n1753) );
  CLKNAND2X2 U1420 ( .A(n1268), .B(n2110), .Y(n412) );
  ADDFX1 U1421 ( .A(n2139), .B(fu_ALU_o1reg[23]), .CI(
        fu_ALU_fu_arch_add_171_carry_23_), .CO(
        fu_ALU_fu_arch_add_171_carry_24_), .S(fu_ALU_fu_arch_N56) );
  ADDFX1 U1422 ( .A(n2162), .B(fu_ALU_o1reg[10]), .CI(
        fu_ALU_fu_arch_add_171_carry_10_), .CO(
        fu_ALU_fu_arch_add_171_carry_11_), .S(fu_ALU_fu_arch_N43) );
  NAND2X2 U1423 ( .A(fu_ALU_fu_arch_n111), .B(fu_ALU_fu_arch_n142), .Y(
        fu_ALU_fu_arch_n141) );
  CLKBUFX4 U1424 ( .A(fu_ALU_fu_arch_n479), .Y(n1829) );
  INVX10 U1425 ( .A(n2127), .Y(fu_ALU_fu_arch_sub_200_B_29_) );
  BUFX18 U1426 ( .A(fu_ALU_fu_arch_n175), .Y(n1762) );
  INVX8 U1427 ( .A(fu_ALU_fu_arch_sub_200_B_27_), .Y(n1764) );
  INVX4 U1428 ( .A(fu_ALU_o1reg[19]), .Y(n2146) );
  BUFX8 U1429 ( .A(rf_RF_t1data_wire[29]), .Y(n1861) );
  OAI211X2 U1430 ( .A0(n1869), .A1(n1764), .B0(fu_ALU_fu_arch_n382), .C0(
        fu_ALU_fu_arch_n383), .Y(ic_socket_ALU_o1_data0_wire[27]) );
  AOI21X1 U1431 ( .A0(n2193), .A1(fu_ALU_fu_arch_N62), .B0(fu_ALU_fu_arch_n354), .Y(fu_ALU_fu_arch_n338) );
  ADDFX1 U1432 ( .A(n2128), .B(n2127), .CI(fu_ALU_fu_arch_sub_200_carry_29_), 
        .CO(fu_ALU_fu_arch_sub_200_carry_30_), .S(fu_ALU_fu_arch_N641) );
  AOI21X1 U1433 ( .A0(n2193), .A1(fu_ALU_fu_arch_N61), .B0(fu_ALU_fu_arch_n374), .Y(fu_ALU_fu_arch_n359) );
  ADDFX1 U1434 ( .A(n2130), .B(n2129), .CI(fu_ALU_fu_arch_sub_200_carry_28_), 
        .CO(fu_ALU_fu_arch_sub_200_carry_29_), .S(fu_ALU_fu_arch_N640) );
  INVX2 U1435 ( .A(n571), .Y(n1894) );
  BUFX8 U1436 ( .A(n219), .Y(n2121) );
  OAI222X1 U1437 ( .A0(fu_ALU_fu_arch_n351), .A1(fu_ALU_fu_arch_n212), .B0(
        fu_ALU_fu_arch_n133), .B1(fu_ALU_fu_arch_n138), .C0(
        fu_ALU_fu_arch_n621), .C1(fu_ALU_fu_arch_n671), .Y(fu_ALU_fu_arch_n659) );
  AOI21X1 U1438 ( .A0(fu_ALU_o1reg[29]), .A1(n2202), .B0(fu_ALU_fu_arch_n312), 
        .Y(fu_ALU_fu_arch_n728) );
  NOR2X5 U1439 ( .A(n2172), .B(n2106), .Y(fu_ALU_fu_arch_n278) );
  NAND2X2 U1440 ( .A(n1779), .B(fu_ALU_fu_arch_sub_200_A_1_), .Y(n2107) );
  NAND2X6 U1441 ( .A(n1779), .B(fu_ALU_fu_arch_sub_200_A_1_), .Y(n2108) );
  INVX4 U1442 ( .A(fu_ALU_fu_arch_sub_200_B_18_), .Y(n1771) );
  NAND2BX2 U1443 ( .AN(n2130), .B(fu_ALU_fu_arch_lt_gt_188_A_28_), .Y(n2019)
         );
  INVX8 U1444 ( .A(n2167), .Y(n1766) );
  INVX6 U1445 ( .A(n2154), .Y(n1767) );
  INVX5 U1446 ( .A(n2173), .Y(n1773) );
  INVX10 U1447 ( .A(n2174), .Y(n1768) );
  INVX5 U1448 ( .A(n2128), .Y(n1765) );
  INVX10 U1449 ( .A(n2171), .Y(fu_ALU_fu_arch_sub_200_B_4_) );
  BUFX10 U1450 ( .A(fu_ALU_o1reg[16]), .Y(n2151) );
  CLKBUFX16 U1451 ( .A(fu_ALU_o1reg[7]), .Y(n2166) );
  INVX4 U1452 ( .A(fu_ALU_o1reg[14]), .Y(n2155) );
  BUFX8 U1453 ( .A(fu_ALU_t1reg[29]), .Y(n2128) );
  BUFX8 U1454 ( .A(fu_ALU_o1reg[27]), .Y(fu_ALU_fu_arch_sub_200_B_27_) );
  ADDFX1 U1455 ( .A(n2128), .B(fu_ALU_o1reg[29]), .CI(
        fu_ALU_fu_arch_add_171_carry_29_), .CO(
        fu_ALU_fu_arch_add_171_carry_30_), .S(fu_ALU_fu_arch_N62) );
  AOI22X2 U1456 ( .A0(n1852), .A1(n1812), .B0(n2121), .B1(
        fu_LSU_o1shadow_reg_9_), .Y(n112) );
  INVX8 U1457 ( .A(n1809), .Y(n1810) );
  INVX12 U1458 ( .A(n2096), .Y(n2110) );
  AND4X2 U1459 ( .A(n378), .B(n379), .C(n380), .D(n381), .Y(n1824) );
  OAI22X1 U1460 ( .A0(fu_ALU_fu_arch_n510), .A1(fu_ALU_fu_arch_n463), .B0(
        fu_ALU_fu_arch_n213), .B1(fu_ALU_fu_arch_n430), .Y(fu_ALU_fu_arch_n509) );
  CLKBUFX4 U1461 ( .A(fu_ALU_fu_arch_n347), .Y(n1882) );
  INVX5 U1462 ( .A(n1833), .Y(fu_ALU_fu_arch_n138) );
  AOI211X2 U1463 ( .A0(n1954), .A1(n1953), .B0(n1952), .C0(n1951), .Y(n2016)
         );
  INVX4 U1464 ( .A(n1776), .Y(fu_ALU_fu_arch_n255) );
  BUFX12 U1465 ( .A(fu_ALU_fu_arch_n281), .Y(n1776) );
  NOR3BX2 U1466 ( .AN(n2137), .B(n2012), .C(n2136), .Y(n1946) );
  OAI21X3 U1467 ( .A0(n1771), .A1(n2149), .B0(n2074), .Y(n2078) );
  OAI21X3 U1468 ( .A0(n1771), .A1(n2149), .B0(n1999), .Y(n2003) );
  CLKBUFX16 U1469 ( .A(fu_ALU_fu_arch_n129), .Y(n2191) );
  NOR3BX2 U1470 ( .AN(n2162), .B(n1978), .C(n2161), .Y(n1979) );
  NOR3BX2 U1471 ( .AN(n2137), .B(n2087), .C(n2136), .Y(n2020) );
  NOR3BX2 U1472 ( .AN(n2152), .B(n2071), .C(n2151), .Y(n2072) );
  NOR3BX2 U1473 ( .AN(n2152), .B(n1997), .C(n2151), .Y(n1998) );
  AND2X4 U1474 ( .A(fu_ALU_fu_arch_sub_200_A_1_), .B(n2184), .Y(n2095) );
  AND2X2 U1475 ( .A(n1779), .B(n2181), .Y(fu_ALU_fu_arch_add_171_carry_1_) );
  INVX14 U1476 ( .A(fu_ALU_fu_arch_sub_200_A_1_), .Y(n1770) );
  INVX2 U1477 ( .A(fu_ALU_fu_arch_sub_200_B_2_), .Y(
        fu_ALU_fu_arch_sub_200_B_not_2_) );
  OR2X2 U1478 ( .A(fu_ALU_fu_arch_sub_200_B_not_0_), .B(n1779), .Y(
        fu_ALU_fu_arch_sub_200_carry_1_) );
  INVX8 U1479 ( .A(n2124), .Y(n1774) );
  INVX4 U1480 ( .A(n2161), .Y(n1772) );
  INVX20 U1481 ( .A(n2178), .Y(fu_ALU_fu_arch_sub_200_A_1_) );
  INVX8 U1482 ( .A(n2148), .Y(fu_ALU_fu_arch_sub_200_B_18_) );
  INVX10 U1483 ( .A(n2142), .Y(fu_ALU_fu_arch_sub_200_B_21_) );
  CLKNAND2X12 U1484 ( .A(inst_fetch_ra_load_wire), .B(n2208), .Y(n264) );
  INVX8 U1485 ( .A(n2132), .Y(n1763) );
  INVX10 U1486 ( .A(fu_ALU_o1reg[13]), .Y(fu_ALU_fu_arch_n621) );
  BUFX8 U1487 ( .A(fu_ALU_o1reg[3]), .Y(n2173) );
  INVX5 U1488 ( .A(fu_ALU_o1reg[21]), .Y(n2142) );
  INVX5 U1489 ( .A(fu_ALU_o1reg[22]), .Y(n2140) );
  BUFX8 U1490 ( .A(rf_RF_t1data_wire[30]), .Y(n1862) );
  OAI211X2 U1491 ( .A0(n2259), .A1(n67), .B0(n68), .C0(n69), .Y(
        rf_RF_t1data_wire[29]) );
  OAI211X2 U1492 ( .A0(n1848), .A1(fu_ALU_fu_arch_n270), .B0(
        fu_ALU_fu_arch_n359), .C0(fu_ALU_fu_arch_n360), .Y(
        ic_socket_ALU_o1_data0_wire[28]) );
  OAI211X2 U1493 ( .A0(n1874), .A1(n1763), .B0(fu_ALU_fu_arch_n403), .C0(
        fu_ALU_fu_arch_n404), .Y(ic_socket_ALU_o1_data0_wire[26]) );
  BUFX3 U1494 ( .A(n233), .Y(n1826) );
  AOI21X4 U1495 ( .A0(n2181), .A1(fu_ALU_fu_arch_n739), .B0(
        fu_ALU_fu_arch_n740), .Y(fu_ALU_fu_arch_n738) );
  AND4X2 U1496 ( .A(n398), .B(n399), .C(n400), .D(n401), .Y(n1809) );
  INVX5 U1497 ( .A(n334), .Y(n1852) );
  NAND4X2 U1498 ( .A(fu_ALU_opc1reg[2]), .B(fu_ALU_fu_arch_n751), .C(
        fu_ALU_fu_arch_N99), .D(fu_ALU_fu_arch_n746), .Y(fu_ALU_fu_arch_n750)
         );
  OAI2B2X1 U1499 ( .A1N(n2166), .A0(fu_ALU_fu_arch_n172), .B0(n1880), .B1(
        fu_ALU_fu_arch_n108), .Y(fu_ALU_fu_arch_n171) );
  OAI2B2X1 U1500 ( .A1N(n2168), .A0(fu_ALU_fu_arch_n186), .B0(
        fu_ALU_fu_arch_n187), .B1(fu_ALU_fu_arch_n108), .Y(fu_ALU_fu_arch_n185) );
  AO22X2 U1501 ( .A0(n1775), .A1(n1829), .B0(fu_ALU_fu_arch_n249), .B1(n1828), 
        .Y(n1879) );
  AOI22X2 U1502 ( .A0(n1775), .A1(n1835), .B0(fu_ALU_fu_arch_n249), .B1(n1831), 
        .Y(fu_ALU_fu_arch_n593) );
  BUFX3 U1503 ( .A(fu_ALU_fu_arch_n193), .Y(n1792) );
  NAND2X4 U1504 ( .A(fu_ALU_fu_arch_n658), .B(n1890), .Y(fu_ALU_fu_arch_n435)
         );
  INVX10 U1505 ( .A(fu_ALU_fu_arch_n235), .Y(fu_ALU_fu_arch_n333) );
  BUFX8 U1506 ( .A(fu_ALU_fu_arch_n168), .Y(n2103) );
  CLKBUFX4 U1507 ( .A(fu_ALU_fu_arch_n461), .Y(n1887) );
  INVX6 U1508 ( .A(n1832), .Y(n1833) );
  NAND2X2 U1509 ( .A(n2198), .B(n1780), .Y(n1889) );
  OAI221X2 U1510 ( .A0(n1768), .A1(n2173), .B0(n1959), .B1(
        fu_ALU_fu_arch_sub_200_B_2_), .C0(n1958), .Y(n1963) );
  OAI221X2 U1511 ( .A0(n1768), .A1(n2173), .B0(n2033), .B1(
        fu_ALU_fu_arch_sub_200_B_2_), .C0(n2032), .Y(n2037) );
  BUFX14 U1512 ( .A(n23), .Y(n2250) );
  CLKBUFX4 U1513 ( .A(n2054), .Y(n1783) );
  INVX14 U1514 ( .A(n419), .Y(n39) );
  CLKNAND2X8 U1515 ( .A(n1850), .B(n2172), .Y(fu_ALU_fu_arch_n388) );
  INVX18 U1516 ( .A(fu_ALU_fu_arch_n250), .Y(n2198) );
  BUFX3 U1517 ( .A(n2009), .Y(n1790) );
  BUFX3 U1518 ( .A(n2084), .Y(n1791) );
  NOR2BX4 U1519 ( .AN(fu_ALU_fu_arch_sub_200_B_11_), .B(n2160), .Y(n1978) );
  INVX10 U1520 ( .A(n2172), .Y(fu_ALU_fu_arch_n220) );
  INVX2 U1521 ( .A(fu_ALU_fu_arch_sub_200_B_4_), .Y(
        fu_ALU_fu_arch_sub_200_B_not_4_) );
  INVX12 U1522 ( .A(n2095), .Y(n1769) );
  BUFX14 U1523 ( .A(n59), .Y(n1777) );
  NAND2BX2 U1524 ( .AN(n2130), .B(fu_ALU_fu_arch_lt_gt_188_A_28_), .Y(n1945)
         );
  BUFX5 U1525 ( .A(fu_ALU_fu_arch_n121), .Y(n2189) );
  NAND2X5 U1526 ( .A(n1779), .B(fu_ALU_fu_arch_sub_200_A_1_), .Y(n2093) );
  NOR2X6 U1527 ( .A(rf_RF_r1opcode_wire[0]), .B(n631), .Y(n59) );
  BUFX16 U1528 ( .A(n498), .Y(n2210) );
  INVX8 U1529 ( .A(n2146), .Y(fu_ALU_fu_arch_sub_200_B_19_) );
  INVX8 U1530 ( .A(fu_ALU_fu_arch_sub_200_B_9_), .Y(n1778) );
  INVX2 U1531 ( .A(n2168), .Y(fu_ALU_fu_arch_sub_200_B_not_6_) );
  INVX12 U1532 ( .A(n2125), .Y(fu_ALU_fu_arch_sub_200_B_30_) );
  BUFX8 U1533 ( .A(fu_ALU_t1reg[15]), .Y(n2154) );
  INVX8 U1534 ( .A(fu_ALU_o1reg[17]), .Y(fu_ALU_fu_arch_n522) );
  BUFX10 U1535 ( .A(fu_ALU_t1reg[19]), .Y(n2147) );
  INVX4 U1536 ( .A(fu_ALU_o1reg[25]), .Y(n2134) );
  BUFX12 U1537 ( .A(fu_ALU_t1reg[3]), .Y(n2174) );
  BUFX12 U1538 ( .A(fu_ALU_t1reg[2]), .Y(n2176) );
  BUFX16 U1539 ( .A(fu_ALU_t1reg[4]), .Y(n2172) );
  NAND3X2 U1540 ( .A(fu_ALU_fu_arch_n263), .B(n1781), .C(fu_ALU_fu_arch_n265), 
        .Y(ic_socket_ALU_o1_data0_wire[31]) );
  INVX4 U1541 ( .A(n583), .Y(n581) );
  BUFX8 U1542 ( .A(n539), .Y(n2112) );
  INVX4 U1543 ( .A(n549), .Y(n550) );
  INVX8 U1544 ( .A(n574), .Y(n2207) );
  NOR2X6 U1545 ( .A(inst_decoder_N232), .B(n538), .Y(n530) );
  NOR2X6 U1546 ( .A(n540), .B(n538), .Y(n549) );
  INVX4 U1547 ( .A(n556), .Y(n1859) );
  NAND2X2 U1548 ( .A(n580), .B(n543), .Y(n574) );
  INVX4 U1549 ( .A(n1856), .Y(n543) );
  NOR3X4 U1550 ( .A(n1856), .B(n580), .C(n579), .Y(n590) );
  INVX4 U1551 ( .A(n1894), .Y(n1856) );
  NAND3X4 U1552 ( .A(inst_decoder_instructionword_wire[4]), .B(n566), .C(n540), 
        .Y(n567) );
  INVX8 U1553 ( .A(rf_RF_t1data_wire[14]), .Y(n263) );
  INVX6 U1554 ( .A(rf_RF_t1data_wire[15]), .Y(n254) );
  INVX8 U1555 ( .A(n1823), .Y(n272) );
  INVX8 U1556 ( .A(rf_RF_t1data_wire[11]), .Y(n297) );
  INVX8 U1557 ( .A(n1820), .Y(n286) );
  NAND2X4 U1558 ( .A(n2117), .B(n1270), .Y(n103) );
  AND2X2 U1559 ( .A(n507), .B(n508), .Y(n1885) );
  INVX8 U1560 ( .A(n1822), .Y(n1823) );
  INVX8 U1561 ( .A(n1819), .Y(n1820) );
  INVX8 U1562 ( .A(n1821), .Y(n365) );
  INVX12 U1563 ( .A(n2111), .Y(n220) );
  INVX8 U1564 ( .A(n1816), .Y(n308) );
  INVX8 U1565 ( .A(n1815), .Y(n1816) );
  INVX8 U1566 ( .A(n1812), .Y(n321) );
  AND2X2 U1567 ( .A(n300), .B(n301), .Y(n1883) );
  INVX8 U1568 ( .A(n1811), .Y(n1812) );
  INVX8 U1569 ( .A(n1808), .Y(n385) );
  INVX8 U1570 ( .A(n1810), .Y(n395) );
  AOI211X2 U1571 ( .A0(fu_LSU_t1opcode_wire[1]), .A1(n2183), .B0(n2117), .C0(
        n2248), .Y(n408) );
  AOI22X2 U1572 ( .A0(n2192), .A1(fu_ALU_fu_arch_N627), .B0(
        fu_ALU_fu_arch_n635), .B1(fu_ALU_fu_arch_n636), .Y(fu_ALU_fu_arch_n634) );
  INVX8 U1573 ( .A(n1825), .Y(n375) );
  INVX8 U1574 ( .A(n1818), .Y(n355) );
  INVX8 U1575 ( .A(n1814), .Y(n345) );
  INVX4 U1576 ( .A(rf_RF_t1data_wire[8]), .Y(n333) );
  INVX8 U1577 ( .A(n1824), .Y(n1825) );
  INVX8 U1578 ( .A(n1813), .Y(n1814) );
  INVX8 U1579 ( .A(n1817), .Y(n1818) );
  BUFX14 U1580 ( .A(n472), .Y(n2119) );
  BUFX14 U1581 ( .A(n31), .Y(n2120) );
  BUFX14 U1582 ( .A(n28), .Y(n2123) );
  INVX8 U1583 ( .A(n1900), .Y(n462) );
  AOI22X2 U1584 ( .A0(fu_ALU_fu_arch_n111), .A1(fu_ALU_fu_arch_n190), .B0(
        fu_ALU_fu_arch_n178), .B1(fu_ALU_fu_arch_n191), .Y(fu_ALU_fu_arch_n182) );
  NAND2X2 U1585 ( .A(n1805), .B(fu_ALU_fu_arch_n500), .Y(fu_ALU_fu_arch_n214)
         );
  AOI22X2 U1586 ( .A0(fu_ALU_fu_arch_n111), .A1(fu_ALU_fu_arch_n177), .B0(
        fu_ALU_fu_arch_n178), .B1(fu_ALU_fu_arch_n179), .Y(fu_ALU_fu_arch_n158) );
  BUFX12 U1587 ( .A(n2248), .Y(n2249) );
  INVX8 U1588 ( .A(n2118), .Y(n453) );
  AOI32X2 U1589 ( .A0(n1881), .A1(n2090), .A2(n2089), .B0(n2088), .B1(n1881), 
        .Y(fu_ALU_fu_arch_N99) );
  NOR2X4 U1590 ( .A(fu_ALU_fu_arch_n762), .B(fu_ALU_fu_arch_n763), .Y(
        fu_ALU_fu_arch_n607) );
  OAI21X4 U1591 ( .A0(fu_ALU_fu_arch_n298), .A1(n2203), .B0(
        fu_ALU_fu_arch_n727), .Y(fu_ALU_fu_arch_n416) );
  INVX2 U1592 ( .A(fu_ALU_fu_arch_n435), .Y(fu_ALU_fu_arch_n519) );
  AOI2BB2X2 U1593 ( .B0(n2103), .B1(n1831), .A0N(fu_ALU_fu_arch_n138), .A1N(
        fu_ALU_fu_arch_n195), .Y(fu_ALU_fu_arch_n180) );
  OR2X2 U1594 ( .A(n1870), .B(n1871), .Y(n1869) );
  OR2X2 U1595 ( .A(n1865), .B(n1866), .Y(n1864) );
  OAI2BB2X2 U1596 ( .B0(fu_ALU_fu_arch_n166), .B1(fu_ALU_fu_arch_n138), .A0N(
        n1839), .A1N(n2103), .Y(fu_ALU_fu_arch_n165) );
  BUFX3 U1597 ( .A(fu_ALU_fu_arch_n346), .Y(n1796) );
  OR2X2 U1598 ( .A(n1875), .B(n1876), .Y(n1874) );
  AOI211X2 U1599 ( .A0(n1806), .A1(n454), .B0(n2212), .C0(n495), .Y(n494) );
  NOR2X2 U1600 ( .A(n2212), .B(n1899), .Y(n1898) );
  BUFX3 U1601 ( .A(fu_ALU_fu_arch_n368), .Y(n1795) );
  BUFX3 U1602 ( .A(fu_ALU_fu_arch_n314), .Y(n1794) );
  NOR2X2 U1603 ( .A(n2190), .B(n1868), .Y(n1866) );
  NOR2X2 U1604 ( .A(n2190), .B(n1873), .Y(n1871) );
  BUFX3 U1605 ( .A(fu_ALU_fu_arch_n482), .Y(n1847) );
  NOR2X2 U1606 ( .A(n2190), .B(n1878), .Y(n1876) );
  OAI211X2 U1607 ( .A0(n2142), .A1(n2199), .B0(fu_ALU_fu_arch_n516), .C0(
        fu_ALU_fu_arch_n517), .Y(fu_ALU_fu_arch_n347) );
  NOR2X2 U1608 ( .A(n2190), .B(n1877), .Y(n1875) );
  BUFX3 U1609 ( .A(fu_ALU_fu_arch_n164), .Y(n1800) );
  AOI21X6 U1610 ( .A0(n2202), .A1(fu_ALU_o1reg[20]), .B0(fu_ALU_fu_arch_n669), 
        .Y(fu_ALU_fu_arch_n131) );
  NOR2X2 U1611 ( .A(n2190), .B(n1867), .Y(n1865) );
  NOR2X2 U1612 ( .A(n2190), .B(n1872), .Y(n1870) );
  BUFX3 U1613 ( .A(fu_ALU_fu_arch_n288), .Y(n1793) );
  BUFX3 U1614 ( .A(fu_ALU_fu_arch_n167), .Y(n1839) );
  INVX4 U1615 ( .A(n1848), .Y(fu_ALU_fu_arch_n456) );
  BUFX3 U1616 ( .A(fu_ALU_fu_arch_n287), .Y(n1799) );
  OAI22X1 U1617 ( .A0(n1848), .A1(fu_ALU_fu_arch_n544), .B0(n1844), .B1(
        fu_ALU_fu_arch_n468), .Y(fu_ALU_fu_arch_n763) );
  BUFX3 U1618 ( .A(fu_ALU_fu_arch_n315), .Y(n1801) );
  AOI21X6 U1619 ( .A0(n2197), .A1(n2157), .B0(fu_ALU_fu_arch_n756), .Y(
        fu_ALU_fu_arch_n155) );
  INVX8 U1620 ( .A(n1853), .Y(n1854) );
  INVX4 U1621 ( .A(n1802), .Y(fu_ALU_fu_arch_n334) );
  OAI22X1 U1622 ( .A0(fu_ALU_fu_arch_n618), .A1(fu_ALU_fu_arch_n617), .B0(
        fu_ALU_fu_arch_n619), .B1(fu_ALU_fu_arch_n563), .Y(fu_ALU_fu_arch_n613) );
  AND2X2 U1623 ( .A(fu_ALU_fu_arch_n350), .B(n1889), .Y(n1890) );
  AOI22X2 U1624 ( .A0(n2202), .A1(fu_ALU_fu_arch_lt_gt_188_A_28_), .B0(n2200), 
        .B1(n2132), .Y(fu_ALU_fu_arch_n658) );
  BUFX14 U1625 ( .A(n19), .Y(n2254) );
  BUFX14 U1626 ( .A(n19), .Y(n2255) );
  CLKBUFX4 U1627 ( .A(fu_ALU_fu_arch_n358), .Y(n1848) );
  NOR2X2 U1628 ( .A(fu_ALU_fu_arch_n544), .B(n1797), .Y(fu_ALU_fu_arch_n168)
         );
  OR2X2 U1629 ( .A(n2133), .B(fu_ALU_fu_arch_n417), .Y(n1877) );
  AOI2BB2X2 U1630 ( .B0(n2057), .B1(n2056), .A0N(n2055), .A1N(n1783), .Y(n2058) );
  OR2X2 U1631 ( .A(n2099), .B(fu_ALU_fu_arch_n417), .Y(n1878) );
  INVX10 U1632 ( .A(fu_ALU_fu_arch_n601), .Y(fu_ALU_fu_arch_n395) );
  AOI2BB2X2 U1633 ( .B0(n1983), .B1(n1982), .A0N(n1981), .A1N(n1784), .Y(n1984) );
  OR2X2 U1634 ( .A(n2131), .B(fu_ALU_fu_arch_n400), .Y(n1872) );
  OR2X2 U1635 ( .A(n2150), .B(fu_ALU_fu_arch_n598), .Y(n1867) );
  OR2X2 U1636 ( .A(n2188), .B(fu_ALU_fu_arch_n598), .Y(n1868) );
  OR2X2 U1637 ( .A(n2188), .B(fu_ALU_fu_arch_n400), .Y(n1873) );
  BUFX14 U1638 ( .A(n276), .Y(n2113) );
  NOR2X2 U1639 ( .A(n521), .B(n2252), .Y(n23) );
  NOR2X6 U1640 ( .A(fu_ALU_fu_arch_n249), .B(n1774), .Y(fu_ALU_fu_arch_n648)
         );
  AND3X2 U1641 ( .A(n1942), .B(n1941), .C(n1940), .Y(fu_ALU_fu_arch_N97) );
  NAND2X4 U1642 ( .A(n2197), .B(n2124), .Y(fu_ALU_fu_arch_n283) );
  CLKBUFX40 U1643 ( .A(fu_ALU_fu_arch_n255), .Y(n2200) );
  BUFX14 U1644 ( .A(n39), .Y(n2246) );
  BUFX8 U1645 ( .A(fu_ALU_fu_arch_n391), .Y(n2100) );
  NOR2X4 U1646 ( .A(n2133), .B(n2195), .Y(fu_ALU_fu_arch_n417) );
  AND2X2 U1647 ( .A(n302), .B(n303), .Y(n1884) );
  NOR2X4 U1648 ( .A(n2131), .B(n2195), .Y(fu_ALU_fu_arch_n400) );
  AOI222X2 U1649 ( .A0(n2197), .A1(fu_ALU_fu_arch_sub_200_B_2_), .B0(n2181), 
        .B1(n2201), .C0(n2177), .C1(fu_ALU_fu_arch_n255), .Y(
        fu_ALU_fu_arch_n580) );
  INVX8 U1650 ( .A(fu_ALU_fu_arch_n430), .Y(fu_ALU_fu_arch_n240) );
  BUFX14 U1651 ( .A(n2242), .Y(n2240) );
  BUFX5 U1652 ( .A(n2188), .Y(n2099) );
  INVX20 U1653 ( .A(n2199), .Y(n2197) );
  BUFX14 U1654 ( .A(n2230), .Y(n2228) );
  INVX2 U1655 ( .A(n2040), .Y(n2043) );
  BUFX14 U1656 ( .A(n2238), .Y(n2237) );
  BUFX14 U1657 ( .A(n2238), .Y(n2236) );
  INVX2 U1658 ( .A(n1966), .Y(n1969) );
  BUFX14 U1659 ( .A(n2226), .Y(n2225) );
  BUFX14 U1660 ( .A(n2242), .Y(n2241) );
  OR2X2 U1661 ( .A(n452), .B(n446), .Y(n1899) );
  BUFX14 U1662 ( .A(n2230), .Y(n2227) );
  BUFX3 U1663 ( .A(n2002), .Y(n1785) );
  BUFX14 U1664 ( .A(n2234), .Y(n2233) );
  BUFX14 U1665 ( .A(n2234), .Y(n2232) );
  BUFX14 U1666 ( .A(n2234), .Y(n2231) );
  BUFX14 U1667 ( .A(n2226), .Y(n2223) );
  BUFX14 U1668 ( .A(n2230), .Y(n2229) );
  BUFX14 U1669 ( .A(n2238), .Y(n2235) );
  BUFX3 U1670 ( .A(n2077), .Y(n1786) );
  BUFX14 U1671 ( .A(n2242), .Y(n2239) );
  BUFX14 U1672 ( .A(n2226), .Y(n2224) );
  AND2X2 U1673 ( .A(n509), .B(n510), .Y(n1886) );
  OAI2B11X2 U1674 ( .A1N(fu_ALU_fu_arch_sub_200_B_29_), .A0(n2128), .B0(n1945), 
        .C0(n1954), .Y(n2009) );
  OAI2B11X2 U1675 ( .A1N(fu_ALU_fu_arch_sub_200_B_21_), .A0(n2143), .B0(n1992), 
        .C0(n2008), .Y(n2002) );
  OAI2B11X2 U1676 ( .A1N(fu_ALU_fu_arch_sub_200_B_21_), .A0(n2143), .B0(n2066), 
        .C0(n2083), .Y(n2077) );
  BUFX14 U1677 ( .A(n47), .Y(n2226) );
  BUFX14 U1678 ( .A(n45), .Y(n2234) );
  BUFX14 U1679 ( .A(n626), .Y(n2205) );
  BUFX14 U1680 ( .A(n626), .Y(n2204) );
  BUFX14 U1681 ( .A(n46), .Y(n2230) );
  BUFX14 U1682 ( .A(n43), .Y(n2242) );
  BUFX14 U1683 ( .A(n44), .Y(n2238) );
  OAI22X1 U1684 ( .A0(n1950), .A1(fu_ALU_fu_arch_sub_200_B_30_), .B0(n1774), 
        .B1(n2180), .Y(n1951) );
  NAND2X4 U1685 ( .A(n2210), .B(n2185), .Y(n419) );
  CLKBUFX16 U1686 ( .A(fu_ALU_fu_arch_n248), .Y(n2104) );
  OAI22X1 U1687 ( .A0(n2004), .A1(fu_ALU_o1reg[22]), .B0(n1737), .B1(n2138), 
        .Y(n2005) );
  OR2X6 U1688 ( .A(fu_ALU_fu_arch_n760), .B(n2189), .Y(n2092) );
  NAND3X2 U1689 ( .A(n1916), .B(n1915), .C(n1914), .Y(n1937) );
  INVX20 U1690 ( .A(n2203), .Y(n1775) );
  OAI2B11X2 U1691 ( .A1N(fu_ALU_fu_arch_sub_200_B_29_), .A0(n2128), .B0(n2019), 
        .C0(n2028), .Y(n2084) );
  INVX6 U1692 ( .A(fu_ALU_fu_arch_n212), .Y(fu_ALU_fu_arch_n111) );
  INVX20 U1693 ( .A(n2189), .Y(n2188) );
  INVX20 U1694 ( .A(n2210), .Y(n2211) );
  INVX8 U1695 ( .A(fu_ALU_fu_arch_n292), .Y(fu_ALU_fu_arch_n242) );
  OAI2B11X2 U1696 ( .A1N(fu_ALU_o1reg[13]), .A0(n2156), .B0(n2047), .C0(n2062), 
        .Y(n2054) );
  CLKAND2X4 U1697 ( .A(n2210), .B(fu_ALU_t1load_wire), .Y(n2098) );
  OAI22X1 U1698 ( .A0(n1974), .A1(n2157), .B0(n1740), .B1(fu_ALU_o1reg[13]), 
        .Y(n1987) );
  BUFX14 U1699 ( .A(n266), .Y(n2115) );
  AO2B2X2 U1700 ( .B0(n2166), .B1(n1766), .A0(fu_ALU_o1reg[6]), .A1N(n2169), 
        .Y(n1968) );
  AO2B2X2 U1701 ( .B0(n2166), .B1(n1766), .A0(n2168), .A1N(n2169), .Y(n2042)
         );
  BUFX12 U1702 ( .A(n2215), .Y(n2216) );
  OA22X2 U1703 ( .A0(n1965), .A1(fu_ALU_fu_arch_sub_200_B_5_), .B0(n1964), 
        .B1(fu_ALU_fu_arch_sub_200_B_4_), .Y(n1970) );
  CLKBUFX6 U1704 ( .A(n2107), .Y(n2109) );
  NAND2X2 U1705 ( .A(inst_fetch_N79), .B(n2208), .Y(n626) );
  OA22X2 U1706 ( .A0(n2039), .A1(fu_ALU_fu_arch_sub_200_B_5_), .B0(n2038), 
        .B1(fu_ALU_o1reg[4]), .Y(n2044) );
  CLKXOR2X2 U1707 ( .A(fu_ALU_fu_arch_sub_200_B_18_), .B(n2149), .Y(n1938) );
  XOR2X1 U1708 ( .A(fu_ALU_o1reg[3]), .B(n2174), .Y(n1908) );
  CLKXOR2X2 U1709 ( .A(fu_ALU_fu_arch_sub_200_B_27_), .B(n2131), .Y(n1918) );
  CLKXOR2X2 U1710 ( .A(n2161), .B(n2162), .Y(n1922) );
  NAND2X2 U1711 ( .A(n2039), .B(fu_ALU_fu_arch_sub_200_B_5_), .Y(n2036) );
  INVX2 U1712 ( .A(fu_ALU_fu_arch_sub_200_B_30_), .Y(
        fu_ALU_fu_arch_sub_200_B_not_30_) );
  OR3X2 U1713 ( .A(fu_ALU_opc1reg[0]), .B(fu_ALU_opc1reg[1]), .C(
        fu_ALU_fu_arch_n745), .Y(fu_ALU_fu_arch_n378) );
  INVX2 U1714 ( .A(n2138), .Y(fu_ALU_fu_arch_sub_200_B_not_23_) );
  INVX2 U1715 ( .A(fu_ALU_fu_arch_sub_200_B_22_), .Y(
        fu_ALU_fu_arch_sub_200_B_not_22_) );
  INVX2 U1716 ( .A(fu_ALU_fu_arch_sub_200_B_21_), .Y(
        fu_ALU_fu_arch_sub_200_B_not_21_) );
  INVX2 U1717 ( .A(n2144), .Y(fu_ALU_fu_arch_sub_200_B_not_20_) );
  INVX2 U1718 ( .A(n2151), .Y(fu_ALU_fu_arch_sub_200_B_not_16_) );
  INVX2 U1719 ( .A(n2157), .Y(fu_ALU_fu_arch_sub_200_B_not_12_) );
  CLKNAND2X2 U1720 ( .A(n1965), .B(fu_ALU_fu_arch_sub_200_B_5_), .Y(n1962) );
  INVX12 U1721 ( .A(n2185), .Y(n132) );
  CLKBUFX16 U1722 ( .A(n58), .Y(n2215) );
  NOR2X2 U1723 ( .A(n586), .B(n585), .Y(n52) );
  OR3X2 U1724 ( .A(fu_ALU_opc1reg[3]), .B(fu_ALU_opc1reg[1]), .C(
        fu_ALU_fu_arch_n746), .Y(fu_ALU_fu_arch_n121) );
  CLKBUFX24 U1725 ( .A(fu_ALU_fu_arch_n130), .Y(n2193) );
  INVX4 U1726 ( .A(n2140), .Y(fu_ALU_fu_arch_sub_200_B_22_) );
  INVX12 U1727 ( .A(n149), .Y(n2187) );
  INVX2 U1728 ( .A(fu_ALU_o1reg[17]), .Y(fu_ALU_fu_arch_sub_200_B_not_17_) );
  BUFX14 U1729 ( .A(ic_socket_gcu_o1_bus_cntrl_wire_0_), .Y(n2186) );
  NAND2X4 U1730 ( .A(inst_decoder_N121), .B(inst_decoder_N230), .Y(n553) );
  INVX4 U1731 ( .A(fu_ALU_t1reg[5]), .Y(n1965) );
  BUFX8 U1732 ( .A(fu_ALU_o1reg[31]), .Y(n2124) );
  BUFX8 U1733 ( .A(fu_ALU_o1reg[6]), .Y(n2168) );
  BUFX8 U1734 ( .A(fu_ALU_t1reg[7]), .Y(n2167) );
  BUFX10 U1735 ( .A(fu_ALU_o1reg[23]), .Y(n2138) );
  INVX10 U1736 ( .A(ic_socket_lsu_o1_bus_cntrl_wire_0_), .Y(n149) );
  BUFX10 U1737 ( .A(fu_ALU_o1reg[12]), .Y(n2157) );
  BUFX10 U1738 ( .A(fu_ALU_t1reg[22]), .Y(n2141) );
  BUFX10 U1739 ( .A(fu_ALU_t1reg[14]), .Y(n2179) );
  BUFX14 U1740 ( .A(fu_ALU_o1reg[15]), .Y(n2153) );
  BUFX10 U1741 ( .A(fu_ALU_o1reg[20]), .Y(n2144) );
  BUFX10 U1742 ( .A(fu_ALU_t1reg[20]), .Y(n2145) );
  BUFX8 U1743 ( .A(fu_ALU_o1reg[10]), .Y(n2161) );
  BUFX10 U1744 ( .A(fu_ALU_t1reg[10]), .Y(n2162) );
  BUFX10 U1745 ( .A(fu_ALU_t1reg[11]), .Y(n2160) );
  BUFX10 U1746 ( .A(fu_ALU_t1reg[16]), .Y(n2152) );
  BUFX10 U1747 ( .A(fu_ALU_t1reg[17]), .Y(n2150) );
  BUFX10 U1748 ( .A(fu_ALU_t1reg[18]), .Y(n2149) );
  INVX4 U1749 ( .A(fu_ALU_o1reg[8]), .Y(n2164) );
  INVX4 U1750 ( .A(fu_ALU_o1reg[29]), .Y(n2127) );
  BUFX10 U1751 ( .A(fu_ALU_t1reg[27]), .Y(n2131) );
  BUFX10 U1752 ( .A(fu_ALU_t1reg[26]), .Y(n2133) );
  BUFX10 U1753 ( .A(fu_ALU_t1reg[30]), .Y(n2126) );
  BUFX8 U1754 ( .A(fu_ALU_o1reg[26]), .Y(n2132) );
  BUFX8 U1755 ( .A(fu_ALU_o1reg[24]), .Y(n2136) );
  BUFX10 U1756 ( .A(fu_ALU_t1reg[25]), .Y(n2135) );
  BUFX10 U1757 ( .A(fu_LSU_o1load_wire), .Y(n2185) );
  BUFX10 U1758 ( .A(fu_ALU_t1reg[24]), .Y(n2137) );
  OR2X2 U1759 ( .A(fu_LSU_status_addr_reg_1__1_), .B(fu_LSU_data_in[23]), .Y(
        n1901) );
  MX2X1 U1760 ( .A(n1808), .B(n2174), .S0(n2252), .Y(n968) );
  MX2X1 U1761 ( .A(n1821), .B(fu_ALU_t1reg[5]), .S0(n2253), .Y(n938) );
  AO21X2 U1762 ( .A0(n1855), .A1(fu_ALU_fu_arch_n249), .B0(fu_ALU_fu_arch_n648), .Y(fu_ALU_fu_arch_n384) );
  INVX5 U1763 ( .A(inst_decoder_N232), .Y(n540) );
  MX2X1 U1764 ( .A(n1825), .B(n2172), .S0(n2252), .Y(n953) );
  OAI2BB1X1 U1765 ( .A0N(fu_LSU_wr_mask_x[7]), .A1N(n2248), .B0(n1274), .Y(
        n1001) );
  OAI2BB1X1 U1766 ( .A0N(fu_LSU_wr_mask_x[30]), .A1N(n2247), .B0(n1278), .Y(
        n1018) );
  OAI2BB1X1 U1767 ( .A0N(fu_LSU_wr_mask_x[5]), .A1N(n2248), .B0(n1274), .Y(
        n1000) );
  OAI2BB1X1 U1768 ( .A0N(fu_LSU_wr_mask_x[28]), .A1N(n2247), .B0(n1278), .Y(
        n1019) );
  OAI2BB1X1 U1769 ( .A0N(fu_LSU_wr_mask_x[3]), .A1N(n2248), .B0(n1274), .Y(
        n999) );
  OAI2BB1X1 U1770 ( .A0N(fu_LSU_wr_mask_x[26]), .A1N(n2247), .B0(n1278), .Y(
        n1020) );
  OAI2BB1X1 U1771 ( .A0N(fu_LSU_wr_mask_x[1]), .A1N(n2248), .B0(n1274), .Y(
        n998) );
  OAI2BB1X1 U1772 ( .A0N(fu_LSU_wr_mask_x[24]), .A1N(n2247), .B0(n1278), .Y(
        n1021) );
  OAI2BB1X1 U1773 ( .A0N(fu_LSU_wr_mask_x[0]), .A1N(n2248), .B0(n1274), .Y(
        n997) );
  OAI2BB1X1 U1774 ( .A0N(fu_LSU_wr_mask_x[25]), .A1N(n2247), .B0(n1278), .Y(
        n1022) );
  OAI2BB1X1 U1775 ( .A0N(fu_LSU_wr_mask_x[2]), .A1N(n2248), .B0(n1274), .Y(
        n996) );
  OAI2BB1X1 U1776 ( .A0N(fu_LSU_wr_mask_x[27]), .A1N(n2247), .B0(n1278), .Y(
        n1023) );
  OAI2BB1X1 U1777 ( .A0N(fu_LSU_wr_mask_x[4]), .A1N(n2248), .B0(n1274), .Y(
        n995) );
  OAI2BB1X1 U1778 ( .A0N(fu_LSU_wr_mask_x[29]), .A1N(n2247), .B0(n1278), .Y(
        n1024) );
  OAI2BB1X1 U1779 ( .A0N(fu_LSU_wr_mask_x[6]), .A1N(n2248), .B0(n1274), .Y(
        n994) );
  OAI2BB1X1 U1780 ( .A0N(fu_LSU_wr_mask_x[31]), .A1N(n2247), .B0(n1278), .Y(
        n1025) );
  OR4X2 U1781 ( .A(n2087), .B(n2086), .C(n2085), .D(n1791), .Y(n2088) );
  OR2X2 U1782 ( .A(n1786), .B(n2078), .Y(n2067) );
  OR2X2 U1783 ( .A(n1785), .B(n2003), .Y(n1993) );
  INVX2 U1784 ( .A(n1783), .Y(n2063) );
  OR4X2 U1785 ( .A(n2012), .B(n2011), .C(n2010), .D(n1790), .Y(n2013) );
  AO22X2 U1786 ( .A0(n1888), .A1(n2101), .B0(n1843), .B1(fu_ALU_fu_arch_n395), 
        .Y(fu_ALU_fu_arch_n585) );
  AO22X2 U1787 ( .A0(n1830), .A1(n2101), .B0(n1828), .B1(fu_ALU_fu_arch_n395), 
        .Y(fu_ALU_fu_arch_n568) );
  AO22X2 U1788 ( .A0(n1849), .A1(fu_ALU_fu_arch_n395), .B0(n1837), .B1(n2101), 
        .Y(fu_ALU_fu_arch_n600) );
  NAND2X2 U1789 ( .A(n1833), .B(fu_ALU_fu_arch_n199), .Y(fu_ALU_fu_arch_n197)
         );
  OR2X2 U1790 ( .A(n2203), .B(n1797), .Y(n1853) );
  OR2X2 U1791 ( .A(n2106), .B(n1797), .Y(n1832) );
  OR2X2 U1792 ( .A(fu_ALU_fu_arch_n468), .B(n1797), .Y(n1891) );
  AOI211X4 U1793 ( .A0(n2083), .A1(n2082), .B0(n2081), .C0(n2080), .Y(n2089)
         );
  CLKXOR2X2 U1794 ( .A(fu_ALU_o1reg[13]), .B(n2156), .Y(n1931) );
  CLKXOR2X2 U1795 ( .A(n2177), .B(fu_ALU_fu_arch_sub_200_A_1_), .Y(n1906) );
  AOI211X4 U1796 ( .A0(n2099), .A1(n2152), .B0(fu_ALU_fu_arch_n620), .C0(n2190), .Y(fu_ALU_fu_arch_n618) );
  CLKXOR2X2 U1797 ( .A(n2151), .B(n2152), .Y(n1902) );
  CLKXOR2X2 U1798 ( .A(fu_ALU_fu_arch_sub_200_B_21_), .B(n2143), .Y(n1907) );
  NOR4X4 U1799 ( .A(fu_ALU_fu_arch_n128), .B(fu_ALU_fu_arch_n678), .C(
        fu_ALU_fu_arch_n679), .D(fu_ALU_fu_arch_n680), .Y(fu_ALU_fu_arch_n677)
         );
  OAI211X2 U1800 ( .A0(n1844), .A1(fu_ALU_fu_arch_n136), .B0(
        fu_ALU_fu_arch_n681), .C0(fu_ALU_fu_arch_n682), .Y(fu_ALU_fu_arch_n680) );
  AOI211X4 U1801 ( .A0(n2104), .A1(fu_ALU_fu_arch_n438), .B0(
        fu_ALU_fu_arch_n518), .C0(fu_ALU_fu_arch_n511), .Y(fu_ALU_fu_arch_n211) );
  NOR2X6 U1802 ( .A(fu_ALU_fu_arch_n544), .B(n1774), .Y(fu_ALU_fu_arch_n518)
         );
  OAI31X4 U1803 ( .A0(n2211), .A1(n605), .A2(n220), .B0(n606), .Y(n1190) );
  XNOR2X2 U1804 ( .A(n1779), .B(fu_ALU_fu_arch_sub_200_B_not_0_), .Y(
        fu_ALU_fu_arch_N612) );
  INVX2 U1805 ( .A(n2181), .Y(fu_ALU_fu_arch_sub_200_B_not_0_) );
  OAI31X4 U1806 ( .A0(inst_decoder_N121), .A1(n537), .A2(n567), .B0(n569), .Y(
        n1145) );
  AOI211X4 U1807 ( .A0(n2169), .A1(fu_ALU_fu_arch_n169), .B0(
        fu_ALU_fu_arch_n184), .C0(fu_ALU_fu_arch_n185), .Y(fu_ALU_fu_arch_n183) );
  AOI211X4 U1808 ( .A0(n2008), .A1(n2007), .B0(n2006), .C0(n2005), .Y(n2014)
         );
  AOI211X4 U1809 ( .A0(n2167), .A1(fu_ALU_fu_arch_n169), .B0(
        fu_ALU_fu_arch_n170), .C0(fu_ALU_fu_arch_n171), .Y(fu_ALU_fu_arch_n159) );
  BUFX2 U1810 ( .A(fu_ALU_fu_arch_n264), .Y(n1781) );
  AOI211X4 U1811 ( .A0(n1775), .A1(fu_ALU_fu_arch_n199), .B0(
        fu_ALU_fu_arch_n542), .C0(fu_ALU_fu_arch_n543), .Y(fu_ALU_fu_arch_n541) );
  CLKXOR2X2 U1812 ( .A(fu_ALU_fu_arch_sub_200_B_2_), .B(n2176), .Y(n1910) );
  CLKXOR2X2 U1813 ( .A(n2166), .B(n2167), .Y(n1927) );
  NAND4X2 U1814 ( .A(n1935), .B(n1934), .C(n1933), .D(n1932), .Y(n1936) );
  NAND4X2 U1815 ( .A(n2269), .B(n2268), .C(n2267), .D(n2266), .Y(n2270) );
  OAI31X4 U1816 ( .A0(fu_LSU_data_in[7]), .A1(n446), .A2(n454), .B0(n496), .Y(
        n495) );
  AOI211X4 U1817 ( .A0(fu_ALU_fu_arch_sub_200_A_1_), .A1(fu_ALU_fu_arch_n169), 
        .B0(fu_ALU_fu_arch_n554), .C0(fu_ALU_fu_arch_n555), .Y(
        fu_ALU_fu_arch_n537) );
  OAI31X4 U1818 ( .A0(n2177), .A1(n1770), .A2(n2195), .B0(fu_ALU_fu_arch_n559), 
        .Y(fu_ALU_fu_arch_n554) );
  NAND4X2 U1819 ( .A(n2265), .B(n2264), .C(n2263), .D(n2262), .Y(n2271) );
  OAI31X4 U1820 ( .A0(n1741), .A1(n2168), .A2(n2195), .B0(fu_ALU_fu_arch_n189), 
        .Y(fu_ALU_fu_arch_n184) );
  AOI22X4 U1821 ( .A0(n2192), .A1(fu_ALU_fu_arch_N617), .B0(n2193), .B1(
        fu_ALU_fu_arch_N38), .Y(fu_ALU_fu_arch_n209) );
  CLKBUFX20 U1822 ( .A(n504), .Y(n2209) );
  CLKXOR2X2 U1823 ( .A(fu_ALU_o1reg[17]), .B(n2150), .Y(n1925) );
  OAI211X2 U1824 ( .A0(fu_ALU_fu_arch_n536), .A1(fu_ALU_fu_arch_n212), .B0(
        fu_ALU_fu_arch_n537), .C0(fu_ALU_fu_arch_n538), .Y(
        ic_socket_ALU_o1_data0_wire[1]) );
  CLKXOR2X2 U1825 ( .A(fu_ALU_fu_arch_sub_200_B_19_), .B(n2147), .Y(n1939) );
  AOI211X4 U1826 ( .A0(n1775), .A1(fu_ALU_fu_arch_n217), .B0(
        fu_ALU_fu_arch_n753), .C0(fu_ALU_fu_arch_n754), .Y(fu_ALU_fu_arch_n741) );
  OAI32X4 U1827 ( .A0(n2106), .A1(n1773), .A2(n2093), .B0(fu_ALU_fu_arch_n757), 
        .B1(n2106), .Y(fu_ALU_fu_arch_n753) );
  CLKXOR2X2 U1828 ( .A(n2132), .B(n2133), .Y(n1911) );
  CLKXOR2X2 U1829 ( .A(fu_ALU_fu_arch_lt_gt_188_A_28_), .B(n2130), .Y(n1919)
         );
  INVX8 U1830 ( .A(n2129), .Y(fu_ALU_fu_arch_lt_gt_188_A_28_) );
  OAI32X4 U1831 ( .A0(fu_ALU_fu_arch_sub_200_B_29_), .A1(n2196), .A2(n1765), 
        .B0(fu_ALU_fu_arch_n356), .B1(n2127), .Y(fu_ALU_fu_arch_n354) );
  BUFX2 U1832 ( .A(n408), .Y(n1782) );
  OAI32X4 U1833 ( .A0(fu_ALU_fu_arch_lt_gt_188_A_28_), .A1(n1747), .A2(n2195), 
        .B0(fu_ALU_fu_arch_n376), .B1(n2129), .Y(fu_ALU_fu_arch_n374) );
  NOR3X6 U1834 ( .A(fu_ALU_fu_arch_n746), .B(fu_ALU_fu_arch_n744), .C(
        fu_ALU_fu_arch_n745), .Y(fu_ALU_fu_arch_n723) );
  INVX2 U1835 ( .A(n1989), .Y(n1784) );
  OAI32X4 U1836 ( .A0(n2003), .A1(n1785), .A2(n2001), .B0(n2000), .B1(n1785), 
        .Y(n2006) );
  OAI32X4 U1837 ( .A0(n2078), .A1(n1786), .A2(n2076), .B0(n2075), .B1(n1786), 
        .Y(n2081) );
  BUFX2 U1838 ( .A(n2016), .Y(n1787) );
  BUFX2 U1839 ( .A(n207), .Y(n1788) );
  NAND4X2 U1840 ( .A(fu_ALU_fu_arch_n715), .B(fu_ALU_fu_arch_n716), .C(
        fu_ALU_fu_arch_n717), .D(fu_ALU_fu_arch_n718), .Y(
        ic_socket_ALU_o1_data0_wire[10]) );
  AOI221X2 U1841 ( .A0(n2162), .A1(fu_ALU_fu_arch_n153), .B0(
        fu_ALU_fu_arch_n719), .B1(fu_ALU_o1reg[10]), .C0(fu_ALU_fu_arch_n720), 
        .Y(fu_ALU_fu_arch_n718) );
  BUFX2 U1842 ( .A(fu_ALU_fu_arch_n211), .Y(n1789) );
  OAI22X2 U1843 ( .A0(n1789), .A1(fu_ALU_fu_arch_n212), .B0(
        fu_ALU_fu_arch_n213), .B1(fu_ALU_fu_arch_n118), .Y(fu_ALU_fu_arch_n201) );
  OAI211X2 U1844 ( .A0(n1789), .A1(fu_ALU_fu_arch_n292), .B0(
        fu_ALU_fu_arch_n503), .C0(fu_ALU_fu_arch_n504), .Y(
        ic_socket_ALU_o1_data0_wire[21]) );
  AOI22X4 U1845 ( .A0(n2198), .A1(fu_ALU_fu_arch_sub_200_B_29_), .B0(n2200), 
        .B1(fu_ALU_fu_arch_sub_200_B_30_), .Y(fu_ALU_fu_arch_n675) );
  OAI211X2 U1846 ( .A0(fu_ALU_fu_arch_n621), .A1(n2108), .B0(
        fu_ALU_fu_arch_n734), .C0(fu_ALU_fu_arch_n735), .Y(fu_ALU_fu_arch_n193) );
  OAI211X2 U1847 ( .A0(n2142), .A1(n1769), .B0(fu_ALU_fu_arch_n466), .C0(
        fu_ALU_fu_arch_n467), .Y(fu_ALU_fu_arch_n288) );
  OAI211X2 U1848 ( .A0(n2140), .A1(n2199), .B0(fu_ALU_fu_arch_n486), .C0(
        fu_ALU_fu_arch_n487), .Y(fu_ALU_fu_arch_n314) );
  OAI211X2 U1849 ( .A0(n2108), .A1(fu_ALU_fu_arch_n522), .B0(
        fu_ALU_fu_arch_n523), .C0(fu_ALU_fu_arch_n524), .Y(fu_ALU_fu_arch_n368) );
  NOR4X4 U1850 ( .A(n1905), .B(n1904), .C(n1903), .D(n1902), .Y(n1942) );
  OAI211X2 U1851 ( .A0(fu_ALU_fu_arch_n522), .A1(n2199), .B0(
        fu_ALU_fu_arch_n604), .C0(fu_ALU_fu_arch_n605), .Y(fu_ALU_fu_arch_n346) );
  NOR4X4 U1852 ( .A(n1909), .B(n1908), .C(n1907), .D(n1906), .Y(n1941) );
  BUFX5 U1853 ( .A(fu_ALU_fu_arch_n608), .Y(n1797) );
  OAI21X1 U1854 ( .A0(fu_ALU_fu_arch_n274), .A1(n1851), .B0(
        fu_ALU_fu_arch_n220), .Y(fu_ALU_fu_arch_n608) );
  CLKBUFX4 U1855 ( .A(fu_ALU_fu_arch_n515), .Y(n1798) );
  AOI22X2 U1856 ( .A0(n2198), .A1(n2177), .B0(n2181), .B1(n2200), .Y(
        fu_ALU_fu_arch_n515) );
  OAI211X2 U1857 ( .A0(fu_ALU_fu_arch_n522), .A1(n1769), .B0(
        fu_ALU_fu_arch_n571), .C0(fu_ALU_fu_arch_n572), .Y(fu_ALU_fu_arch_n287) );
  OAI211X2 U1858 ( .A0(fu_ALU_fu_arch_n621), .A1(n1769), .B0(
        fu_ALU_fu_arch_n705), .C0(fu_ALU_fu_arch_n706), .Y(fu_ALU_fu_arch_n164) );
  OAI211X2 U1859 ( .A0(fu_ALU_fu_arch_n522), .A1(n1776), .B0(
        fu_ALU_fu_arch_n588), .C0(fu_ALU_fu_arch_n589), .Y(fu_ALU_fu_arch_n315) );
  OAI31X4 U1860 ( .A0(inst_decoder_N121), .A1(inst_decoder_N230), .A2(n567), 
        .B0(n570), .Y(n1146) );
  OAI31X4 U1861 ( .A0(fu_LSU_o1load_wire), .A1(n231), .A2(n320), .B0(n331), 
        .Y(n889) );
  AOI211X4 U1862 ( .A0(n132), .A1(n115), .B0(n2182), .C0(n2248), .Y(n416) );
  CLKBUFX4 U1863 ( .A(fu_ALU_fu_arch_n580), .Y(n1802) );
  OAI31X4 U1864 ( .A0(fu_LSU_o1load_wire), .A1(n115), .A2(n103), .B0(n116), 
        .Y(n114) );
  INVX2 U1865 ( .A(fu_ALU_fu_arch_n154), .Y(n1803) );
  INVX4 U1866 ( .A(fu_ALU_fu_arch_n224), .Y(fu_ALU_fu_arch_n154) );
  NOR3X4 U1867 ( .A(rf_RF_r1opcode_wire[1]), .B(n586), .C(n584), .Y(n58) );
  BUFX2 U1868 ( .A(fu_ALU_fu_arch_n262), .Y(n1804) );
  OAI211X2 U1869 ( .A0(n1804), .A1(fu_ALU_fu_arch_n292), .B0(
        fu_ALU_fu_arch_n560), .C0(fu_ALU_fu_arch_n561), .Y(
        ic_socket_ALU_o1_data0_wire[19]) );
  NOR2X4 U1870 ( .A(n1804), .B(fu_ALU_fu_arch_n212), .Y(fu_ALU_fu_arch_n241)
         );
  CLKBUFX4 U1871 ( .A(fu_ALU_fu_arch_n227), .Y(n1805) );
  OAI211X2 U1872 ( .A0(n1805), .A1(fu_ALU_fu_arch_n430), .B0(
        fu_ALU_fu_arch_n520), .C0(fu_ALU_fu_arch_n521), .Y(
        ic_socket_ALU_o1_data0_wire[20]) );
  AOI222X2 U1873 ( .A0(fu_ALU_fu_arch_n457), .A1(n1775), .B0(
        fu_ALU_fu_arch_n534), .B1(fu_ALU_fu_arch_n249), .C0(
        fu_ALU_fu_arch_n456), .C1(n2104), .Y(fu_ALU_fu_arch_n227) );
  CLKBUFX20 U1874 ( .A(n2218), .Y(n2217) );
  CLKBUFX4 U1875 ( .A(n449), .Y(n1806) );
  AOI22X2 U1876 ( .A0(fu_LSU_status_addr_reg_1__1_), .A1(fu_LSU_data_in[15]), 
        .B0(fu_LSU_data_in[31]), .B1(n446), .Y(n449) );
  OAI31X4 U1877 ( .A0(n2196), .A1(n2153), .A2(n1767), .B0(fu_ALU_fu_arch_n634), 
        .Y(fu_ALU_fu_arch_n627) );
  INVX2 U1878 ( .A(fu_ALU_fu_arch_n590), .Y(n1807) );
  OAI211X2 U1879 ( .A0(fu_ALU_fu_arch_n298), .A1(fu_ALU_fu_arch_n270), .B0(
        fu_ALU_fu_arch_n299), .C0(fu_ALU_fu_arch_n300), .Y(fu_ALU_fu_arch_n297) );
  INVX4 U1880 ( .A(fu_ALU_fu_arch_n298), .Y(fu_ALU_fu_arch_n590) );
  AOI211X4 U1881 ( .A0(fu_ALU_fu_arch_lt_gt_188_A_28_), .A1(n2198), .B0(
        fu_ALU_fu_arch_n309), .C0(fu_ALU_fu_arch_n765), .Y(fu_ALU_fu_arch_n358) );
  NOR2X4 U1882 ( .A(n1776), .B(n2127), .Y(fu_ALU_fu_arch_n309) );
  NOR4X4 U1883 ( .A(fu_ALU_fu_arch_n309), .B(fu_ALU_fu_arch_n310), .C(
        fu_ALU_fu_arch_n311), .D(fu_ALU_fu_arch_n312), .Y(fu_ALU_fu_arch_n307)
         );
  NOR2X4 U1884 ( .A(n1769), .B(n2129), .Y(fu_ALU_fu_arch_n312) );
  AOI211X4 U1885 ( .A0(n2177), .A1(n2200), .B0(fu_ALU_fu_arch_n459), .C0(
        fu_ALU_fu_arch_n690), .Y(fu_ALU_fu_arch_n757) );
  AOI211X4 U1886 ( .A0(n2198), .A1(fu_ALU_fu_arch_sub_200_B_4_), .B0(
        fu_ALU_fu_arch_n690), .C0(fu_ALU_fu_arch_n691), .Y(fu_ALU_fu_arch_n461) );
  NOR2X4 U1887 ( .A(n1769), .B(n2175), .Y(fu_ALU_fu_arch_n690) );
  NOR2BX4 U1888 ( .AN(fu_ALU_o1reg[17]), .B(n2150), .Y(n1997) );
  NOR2BX4 U1889 ( .AN(fu_ALU_o1reg[17]), .B(n2150), .Y(n2071) );
  AOI22X2 U1890 ( .A0(n2193), .A1(fu_ALU_fu_arch_N60), .B0(fu_ALU_fu_arch_n399), .B1(fu_ALU_fu_arch_n240), .Y(fu_ALU_fu_arch_n398) );
  NOR2X4 U1891 ( .A(n2174), .B(fu_ALU_fu_arch_n573), .Y(fu_ALU_fu_arch_n399)
         );
  AOI21X4 U1892 ( .A0(fu_LSU_data_out[0]), .A1(n2249), .B0(n413), .Y(n411) );
  OAI32X4 U1893 ( .A0(n250), .A1(n220), .A2(n334), .B0(n235), .B1(n250), .Y(
        n413) );
  AOI21X4 U1894 ( .A0(n2200), .A1(fu_ALU_fu_arch_sub_200_B_8_), .B0(
        fu_ALU_fu_arch_n256), .Y(fu_ALU_fu_arch_n166) );
  OAI211X2 U1895 ( .A0(n1772), .A1(n2109), .B0(fu_ALU_fu_arch_n259), .C0(
        fu_ALU_fu_arch_n260), .Y(fu_ALU_fu_arch_n256) );
  INVX10 U1896 ( .A(n426), .Y(n2213) );
  OAI31X4 U1897 ( .A0(fu_LSU_status_addr_reg_1__3_), .A1(
        fu_LSU_status_addr_reg_1__4_), .A2(fu_LSU_status_addr_reg_1__2_), .B0(
        n497), .Y(n426) );
  OAI32X4 U1898 ( .A0(n2011), .A1(n1790), .A2(n1949), .B0(n1948), .B1(n1790), 
        .Y(n1952) );
  OAI21X4 U1899 ( .A0(n1763), .A1(n2133), .B0(n1947), .Y(n2011) );
  OAI32X4 U1900 ( .A0(n2086), .A1(n1791), .A2(n2023), .B0(n2022), .B1(n1791), 
        .Y(n2026) );
  OAI21X4 U1901 ( .A0(n1763), .A1(n2133), .B0(n2021), .Y(n2086) );
  NOR2BX4 U1902 ( .AN(fu_ALU_fu_arch_sub_200_B_11_), .B(n2160), .Y(n2052) );
  OAI2BB2X4 U1903 ( .B0(n2122), .B1(n334), .A0N(n2121), .A1N(
        fu_LSU_o1shadow_reg_8_), .Y(n129) );
  AOI21X4 U1904 ( .A0(n459), .A1(fu_LSU_status_addr_reg_1__3_), .B0(n457), .Y(
        n470) );
  NOR2BX8 U1905 ( .AN(fu_LSU_status_addr_reg_1__4_), .B(n459), .Y(n457) );
  AOI21X4 U1906 ( .A0(fu_ALU_fu_arch_n249), .A1(fu_ALU_fu_arch_n592), .B0(
        fu_ALU_fu_arch_n648), .Y(fu_ALU_fu_arch_n291) );
  AOI21X4 U1907 ( .A0(fu_ALU_fu_arch_n249), .A1(fu_ALU_fu_arch_n438), .B0(
        fu_ALU_fu_arch_n648), .Y(fu_ALU_fu_arch_n351) );
  OAI211X4 U1908 ( .A0(n2108), .A1(n2142), .B0(fu_ALU_fu_arch_n445), .C0(
        fu_ALU_fu_arch_n446), .Y(fu_ALU_fu_arch_n366) );
  OAI211X4 U1909 ( .A0(n2140), .A1(n2109), .B0(fu_ALU_fu_arch_n421), .C0(
        fu_ALU_fu_arch_n422), .Y(fu_ALU_fu_arch_n345) );
  OAI211X4 U1910 ( .A0(n1763), .A1(n2199), .B0(fu_ALU_fu_arch_n411), .C0(
        fu_ALU_fu_arch_n412), .Y(fu_ALU_fu_arch_n313) );
  OAI211X4 U1911 ( .A0(n1764), .A1(n2199), .B0(fu_ALU_fu_arch_n392), .C0(
        fu_ALU_fu_arch_n393), .Y(fu_ALU_fu_arch_n285) );
  AOI22X2 U1912 ( .A0(n2193), .A1(fu_ALU_fu_arch_N59), .B0(fu_ALU_fu_arch_n240), .B1(fu_ALU_fu_arch_n416), .Y(fu_ALU_fu_arch_n415) );
  OAI211X4 U1913 ( .A0(n1802), .A1(fu_ALU_fu_arch_n544), .B0(
        fu_ALU_fu_arch_n652), .C0(fu_ALU_fu_arch_n653), .Y(fu_ALU_fu_arch_n304) );
  NAND2X2 U1914 ( .A(n2104), .B(n1843), .Y(fu_ALU_fu_arch_n653) );
  NOR4X4 U1915 ( .A(rf_RF_t1opcode_wire[2]), .B(rf_RF_t1opcode_wire[1]), .C(
        n546), .D(n545), .Y(n44) );
  NAND2X5 U1916 ( .A(n2210), .B(rf_RF_t1load_wire), .Y(n545) );
  NOR4X4 U1917 ( .A(rf_RF_t1opcode_wire[2]), .B(n546), .C(n547), .D(n545), .Y(
        n46) );
  CLKBUFX4 U1918 ( .A(rf_RF_t1data_wire[3]), .Y(n1808) );
  NAND4X6 U1919 ( .A(n388), .B(n389), .C(n390), .D(n391), .Y(
        rf_RF_t1data_wire[3]) );
  AND4X2 U1920 ( .A(n324), .B(n325), .C(n326), .D(n327), .Y(n1811) );
  AND4X2 U1921 ( .A(n348), .B(n349), .C(n350), .D(n351), .Y(n1813) );
  AND4X2 U1922 ( .A(n311), .B(n312), .C(n313), .D(n314), .Y(n1815) );
  AND4X2 U1923 ( .A(n358), .B(n359), .C(n360), .D(n361), .Y(n1817) );
  AND4X2 U1924 ( .A(n289), .B(n290), .C(n291), .D(n292), .Y(n1819) );
  CLKBUFX4 U1925 ( .A(rf_RF_t1data_wire[5]), .Y(n1821) );
  NAND4X6 U1926 ( .A(n368), .B(n369), .C(n370), .D(n371), .Y(
        rf_RF_t1data_wire[5]) );
  AND4X2 U1927 ( .A(n278), .B(n279), .C(n280), .D(n281), .Y(n1822) );
  AOI221X4 U1928 ( .A0(fu_LSU_status_addr_reg_1__3_), .A1(
        fu_LSU_status_addr_reg_1__2_), .B0(n458), .B1(n459), .C0(
        fu_LSU_status_addr_reg_1__4_), .Y(n455) );
  NOR4X8 U1929 ( .A(n455), .B(fu_LSU_status_addr_reg_1__0_), .C(n457), .D(
        n2212), .Y(n448) );
  CLKBUFX4 U1930 ( .A(fu_ALU_fu_arch_n192), .Y(n1827) );
  OAI211X2 U1931 ( .A0(fu_ALU_fu_arch_n522), .A1(n2109), .B0(
        fu_ALU_fu_arch_n730), .C0(fu_ALU_fu_arch_n731), .Y(fu_ALU_fu_arch_n192) );
  CLKBUFX4 U1932 ( .A(fu_ALU_fu_arch_n480), .Y(n1828) );
  OAI211X2 U1933 ( .A0(n1754), .A1(n1769), .B0(fu_ALU_fu_arch_n703), .C0(
        fu_ALU_fu_arch_n259), .Y(fu_ALU_fu_arch_n480) );
  OAI211X2 U1934 ( .A0(n1769), .A1(n1738), .B0(fu_ALU_fu_arch_n701), .C0(
        fu_ALU_fu_arch_n551), .Y(fu_ALU_fu_arch_n479) );
  CLKBUFX4 U1935 ( .A(fu_ALU_fu_arch_n474), .Y(n1830) );
  AOI222X4 U1936 ( .A0(n1828), .A1(n1775), .B0(n1830), .B1(fu_ALU_fu_arch_n249), .C0(n1829), .C1(n2104), .Y(fu_ALU_fu_arch_n387) );
  OAI211X2 U1937 ( .A0(n1778), .A1(n1769), .B0(fu_ALU_fu_arch_n702), .C0(
        fu_ALU_fu_arch_n547), .Y(fu_ALU_fu_arch_n474) );
  CLKBUFX4 U1938 ( .A(fu_ALU_fu_arch_n194), .Y(n1831) );
  OAI211X2 U1939 ( .A0(n2142), .A1(n2093), .B0(fu_ALU_fu_arch_n732), .C0(
        fu_ALU_fu_arch_n733), .Y(fu_ALU_fu_arch_n194) );
  AOI211X4 U1940 ( .A0(n1833), .A1(fu_ALU_fu_arch_n217), .B0(
        fu_ALU_fu_arch_n218), .C0(fu_ALU_fu_arch_n219), .Y(fu_ALU_fu_arch_n216) );
  CLKBUFX4 U1941 ( .A(fu_ALU_fu_arch_n162), .Y(n1834) );
  OAI211X2 U1942 ( .A0(fu_ALU_fu_arch_n522), .A1(n1769), .B0(
        fu_ALU_fu_arch_n709), .C0(fu_ALU_fu_arch_n710), .Y(fu_ALU_fu_arch_n162) );
  CLKBUFX4 U1943 ( .A(fu_ALU_fu_arch_n502), .Y(n1835) );
  OAI211X2 U1944 ( .A0(n2140), .A1(n2199), .B0(fu_ALU_fu_arch_n736), .C0(
        fu_ALU_fu_arch_n371), .Y(fu_ALU_fu_arch_n502) );
  CLKBUFX4 U1945 ( .A(fu_ALU_fu_arch_n501), .Y(n1836) );
  AOI22X4 U1946 ( .A0(n1775), .A1(n1836), .B0(fu_ALU_fu_arch_n249), .B1(n1835), 
        .Y(fu_ALU_fu_arch_n488) );
  OAI2BB1X2 U1947 ( .A0N(n2104), .A1N(n1836), .B0(fu_ALU_fu_arch_n593), .Y(
        fu_ALU_fu_arch_n591) );
  OAI211X2 U1948 ( .A0(n1764), .A1(n1776), .B0(fu_ALU_fu_arch_n728), .C0(
        fu_ALU_fu_arch_n729), .Y(fu_ALU_fu_arch_n501) );
  CLKBUFX4 U1949 ( .A(fu_ALU_fu_arch_n440), .Y(n1837) );
  OAI211X2 U1950 ( .A0(n1778), .A1(n2199), .B0(fu_ALU_fu_arch_n667), .C0(
        fu_ALU_fu_arch_n253), .Y(fu_ALU_fu_arch_n440) );
  CLKBUFX4 U1951 ( .A(fu_ALU_fu_arch_n451), .Y(n1838) );
  OAI2BB2X2 U1952 ( .B0(n1887), .B1(fu_ALU_fu_arch_n601), .A0N(n1838), .A1N(
        n2100), .Y(fu_ALU_fu_arch_n611) );
  OAI211X2 U1953 ( .A0(n2108), .A1(n1778), .B0(fu_ALU_fu_arch_n686), .C0(
        fu_ALU_fu_arch_n687), .Y(fu_ALU_fu_arch_n451) );
  CLKBUFX4 U1954 ( .A(fu_ALU_fu_arch_n367), .Y(n1840) );
  OAI211X2 U1955 ( .A0(n2109), .A1(fu_ALU_fu_arch_n621), .B0(
        fu_ALU_fu_arch_n622), .C0(fu_ALU_fu_arch_n623), .Y(fu_ALU_fu_arch_n367) );
  CLKBUFX4 U1956 ( .A(fu_ALU_fu_arch_n396), .Y(n1841) );
  OAI211X2 U1957 ( .A0(fu_ALU_fu_arch_n621), .A1(n1769), .B0(
        fu_ALU_fu_arch_n639), .C0(fu_ALU_fu_arch_n548), .Y(fu_ALU_fu_arch_n396) );
  CLKBUFX4 U1958 ( .A(fu_ALU_fu_arch_n413), .Y(n1842) );
  OAI211X2 U1959 ( .A0(fu_ALU_fu_arch_n621), .A1(n1776), .B0(
        fu_ALU_fu_arch_n654), .C0(fu_ALU_fu_arch_n655), .Y(fu_ALU_fu_arch_n413) );
  CLKBUFX4 U1960 ( .A(fu_ALU_fu_arch_n498), .Y(n1843) );
  AOI22X4 U1961 ( .A0(n1775), .A1(fu_ALU_fu_arch_n334), .B0(
        fu_ALU_fu_arch_n249), .B1(n1843), .Y(fu_ALU_fu_arch_n187) );
  OAI211X2 U1962 ( .A0(n1773), .A1(n2108), .B0(fu_ALU_fu_arch_n725), .C0(
        fu_ALU_fu_arch_n326), .Y(fu_ALU_fu_arch_n498) );
  CLKBUFX4 U1963 ( .A(fu_ALU_fu_arch_n535), .Y(n1844) );
  CLKBUFX4 U1964 ( .A(fu_ALU_fu_arch_n428), .Y(n1845) );
  OAI211X2 U1965 ( .A0(fu_ALU_fu_arch_n621), .A1(n2199), .B0(
        fu_ALU_fu_arch_n666), .C0(fu_ALU_fu_arch_n546), .Y(fu_ALU_fu_arch_n428) );
  CLKBUFX4 U1966 ( .A(fu_ALU_fu_arch_n458), .Y(n1846) );
  AOI222X4 U1967 ( .A0(fu_ALU_fu_arch_n533), .A1(n2174), .B0(n1846), .B1(n1775), .C0(n1838), .C1(fu_ALU_fu_arch_n249), .Y(fu_ALU_fu_arch_n364) );
  OAI211X2 U1968 ( .A0(n1754), .A1(n2108), .B0(fu_ALU_fu_arch_n688), .C0(
        fu_ALU_fu_arch_n689), .Y(fu_ALU_fu_arch_n458) );
  CLKBUFX4 U1969 ( .A(fu_ALU_fu_arch_n439), .Y(n1849) );
  AOI21X4 U1970 ( .A0(n2104), .A1(n1849), .B0(fu_ALU_fu_arch_n664), .Y(
        fu_ALU_fu_arch_n343) );
  OAI211X2 U1971 ( .A0(n2175), .A1(n2093), .B0(fu_ALU_fu_arch_n668), .C0(
        fu_ALU_fu_arch_n550), .Y(fu_ALU_fu_arch_n439) );
  NOR2X2 U1972 ( .A(fu_ALU_opc1reg[0]), .B(fu_ALU_fu_arch_n761), .Y(
        fu_ALU_fu_arch_n266) );
  INVX5 U1973 ( .A(fu_ALU_fu_arch_n378), .Y(n1851) );
  AOI22X4 U1974 ( .A0(n253), .A1(n1816), .B0(n2121), .B1(
        fu_LSU_o1shadow_reg_10_), .Y(n99) );
  AOI22X4 U1975 ( .A0(n1852), .A1(rf_RF_t1data_wire[15]), .B0(n2121), .B1(
        fu_LSU_o1shadow_reg_15_), .Y(n24) );
  AOI22X4 U1976 ( .A0(n1852), .A1(n1820), .B0(n2121), .B1(
        fu_LSU_o1shadow_reg_12_), .Y(n75) );
  AOI22X4 U1977 ( .A0(n1852), .A1(rf_RF_t1data_wire[11]), .B0(n2121), .B1(
        fu_LSU_o1shadow_reg_11_), .Y(n87) );
  AOI22X4 U1978 ( .A0(n1852), .A1(rf_RF_t1data_wire[14]), .B0(n2121), .B1(
        fu_LSU_o1shadow_reg_14_), .Y(n35) );
  AOI22X4 U1979 ( .A0(n1852), .A1(n1823), .B0(n2121), .B1(
        fu_LSU_o1shadow_reg_13_), .Y(n62) );
  INVX4 U1980 ( .A(n253), .Y(n334) );
  NOR2X4 U1981 ( .A(n132), .B(n2249), .Y(n253) );
  INVX4 U1982 ( .A(n1854), .Y(fu_ALU_fu_arch_n134) );
  CLKBUFX4 U1983 ( .A(fu_ALU_fu_arch_n481), .Y(n1855) );
  AOI22X4 U1984 ( .A0(n2176), .A1(fu_ALU_fu_arch_n635), .B0(n1855), .B1(
        fu_ALU_fu_arch_n335), .Y(fu_ALU_fu_arch_n573) );
  AOI22X4 U1985 ( .A0(n1775), .A1(n1855), .B0(fu_ALU_fu_arch_n249), .B1(n1847), 
        .Y(fu_ALU_fu_arch_n469) );
  NOR2X4 U1986 ( .A(n571), .B(n551), .Y(n566) );
  CLKBUFX6 U1987 ( .A(n562), .Y(n1857) );
  NOR2X2 U1988 ( .A(inst_decoder_N232), .B(n552), .Y(n562) );
  CLKBUFX6 U1989 ( .A(n424), .Y(n1858) );
  NOR2X2 U1990 ( .A(n446), .B(n447), .Y(n424) );
  INVX4 U1991 ( .A(n554), .Y(n556) );
  NOR3X6 U1992 ( .A(inst_decoder_N230), .B(n552), .C(n540), .Y(n554) );
  BUFX8 U1993 ( .A(rf_RF_t1data_wire[31]), .Y(n1860) );
  OAI211X2 U1994 ( .A0(n1750), .A1(n513), .B0(n514), .C0(n515), .Y(
        rf_RF_t1data_wire[31]) );
  OAI211X2 U1995 ( .A0(n1750), .A1(n49), .B0(n50), .C0(n51), .Y(
        rf_RF_t1data_wire[30]) );
  OAI31X4 U1996 ( .A0(n2196), .A1(fu_ALU_o1reg[3]), .A2(n1768), .B0(
        fu_ALU_fu_arch_n239), .Y(fu_ALU_fu_arch_n232) );
  OAI31X4 U1997 ( .A0(n2196), .A1(fu_ALU_o1reg[4]), .A2(fu_ALU_fu_arch_n220), 
        .B0(fu_ALU_fu_arch_n223), .Y(fu_ALU_fu_arch_n218) );
  OAI31X4 U1998 ( .A0(n2196), .A1(fu_ALU_o1reg[2]), .A2(fu_ALU_fu_arch_n335), 
        .B0(fu_ALU_fu_arch_n336), .Y(fu_ALU_fu_arch_n329) );
  OAI31X4 U1999 ( .A0(n2196), .A1(n2166), .A2(n1766), .B0(fu_ALU_fu_arch_n176), 
        .Y(fu_ALU_fu_arch_n170) );
  OAI211X2 U2000 ( .A0(n2160), .A1(n2196), .B0(fu_ALU_fu_arch_n704), .C0(n2092), .Y(fu_ALU_fu_arch_n696) );
  INVX12 U2001 ( .A(n1762), .Y(n2196) );
  INVX4 U2002 ( .A(n530), .Y(n532) );
  OAI31X4 U2003 ( .A0(n2110), .A1(n230), .A2(n231), .B0(n232), .Y(n791) );
  INVX2 U2004 ( .A(n1268), .Y(n230) );
  AOI222X4 U2005 ( .A0(n1846), .A1(fu_ALU_fu_arch_n249), .B0(n2104), .B1(
        fu_ALU_fu_arch_n459), .C0(fu_ALU_fu_arch_n460), .C1(n1775), .Y(
        fu_ALU_fu_arch_n139) );
  INVX2 U2006 ( .A(n1887), .Y(fu_ALU_fu_arch_n460) );
  INVX8 U2007 ( .A(n1891), .Y(n1892) );
  NAND2X4 U2008 ( .A(n2174), .B(n2124), .Y(fu_ALU_fu_arch_n437) );
  INVX8 U2009 ( .A(inst_decoder_N121), .Y(n531) );
  OAI22X4 U2010 ( .A0(n2034), .A1(n2168), .B0(n1766), .B1(n2166), .Y(n2040) );
  NOR2X2 U2011 ( .A(n2211), .B(n524), .Y(n276) );
  OAI32X4 U2012 ( .A0(n2211), .A1(n524), .A2(n417), .B0(fu_LSU_wr_en_x[0]), 
        .B1(n2210), .Y(n523) );
  INVX4 U2013 ( .A(fu_LSU_data_in[27]), .Y(n434) );
  INVX4 U2014 ( .A(fu_LSU_data_in[28]), .Y(n437) );
  INVX4 U2015 ( .A(fu_LSU_data_in[26]), .Y(n431) );
  INVX4 U2016 ( .A(fu_LSU_data_in[29]), .Y(n440) );
  INVX4 U2017 ( .A(fu_LSU_data_in[25]), .Y(n428) );
  INVX4 U2018 ( .A(fu_LSU_data_in[30]), .Y(n443) );
  INVX4 U2019 ( .A(fu_LSU_data_in[24]), .Y(n421) );
  NOR3X4 U2020 ( .A(inst_decoder_instructionword_wire[5]), .B(
        inst_decoder_instructionword_wire[4]), .C(n541), .Y(n539) );
  BUFX8 U2021 ( .A(n333), .Y(n2122) );
  AND4X4 U2022 ( .A(fu_ALU_fu_arch_n545), .B(fu_ALU_fu_arch_n546), .C(
        fu_ALU_fu_arch_n547), .D(fu_ALU_fu_arch_n548), .Y(fu_ALU_fu_arch_n137)
         );
  NAND2X2 U2023 ( .A(n2202), .B(n2157), .Y(fu_ALU_fu_arch_n548) );
  NOR4X4 U2024 ( .A(n2185), .B(n239), .C(n2182), .D(n2249), .Y(n31) );
  INVX4 U2025 ( .A(fu_LSU_o1shadow_reg_1_), .Y(n115) );
  INVX4 U2026 ( .A(fu_LSU_o1shadow_reg_0_), .Y(n231) );
  OAI211X2 U2027 ( .A0(fu_ALU_fu_arch_sub_200_B_not_30_), .A1(n1776), .B0(
        fu_ALU_fu_arch_n282), .C0(fu_ALU_fu_arch_n283), .Y(fu_ALU_fu_arch_n279) );
  BUFX2 U2028 ( .A(n2091), .Y(n1881) );
  INVX4 U2029 ( .A(rf_RF_r1opcode_wire[0]), .Y(n584) );
  NOR4X8 U2030 ( .A(rf_RF_r1opcode_wire[0]), .B(rf_RF_r1opcode_wire[1]), .C(
        rf_RF_r1opcode_wire[2]), .D(n1748), .Y(n53) );
  BUFX12 U2031 ( .A(fu_ALU_fu_arch_n247), .Y(n2105) );
  AOI211X4 U2032 ( .A0(n2101), .A1(n1846), .B0(fu_ALU_fu_arch_n296), .C0(
        fu_ALU_fu_arch_n611), .Y(fu_ALU_fu_arch_n610) );
  AOI211X4 U2033 ( .A0(n2100), .A1(n1845), .B0(fu_ALU_fu_arch_n296), .C0(
        fu_ALU_fu_arch_n596), .Y(fu_ALU_fu_arch_n595) );
  AOI211X4 U2034 ( .A0(n2100), .A1(n1842), .B0(fu_ALU_fu_arch_n296), .C0(
        fu_ALU_fu_arch_n579), .Y(fu_ALU_fu_arch_n578) );
  AOI211X4 U2035 ( .A0(n2100), .A1(n1841), .B0(fu_ALU_fu_arch_n296), .C0(
        fu_ALU_fu_arch_n562), .Y(fu_ALU_fu_arch_n561) );
  AOI211X4 U2036 ( .A0(n2101), .A1(n1845), .B0(fu_ALU_fu_arch_n296), .C0(
        fu_ALU_fu_arch_n505), .Y(fu_ALU_fu_arch_n504) );
  INVX8 U2037 ( .A(n2102), .Y(fu_ALU_fu_arch_n296) );
  OAI2BB1X1 U2038 ( .A0N(fu_LSU_wr_mask_x[16]), .A1N(n2247), .B0(n1276), .Y(
        n1013) );
  OAI2BB1X1 U2039 ( .A0N(fu_LSU_wr_mask_x[15]), .A1N(n2248), .B0(n1272), .Y(
        n1009) );
  OAI2BB1X1 U2040 ( .A0N(fu_LSU_wr_mask_x[17]), .A1N(n2247), .B0(n1276), .Y(
        n1014) );
  OAI2BB1X1 U2041 ( .A0N(fu_LSU_wr_mask_x[14]), .A1N(n2248), .B0(n1272), .Y(
        n1002) );
  OAI2BB1X1 U2042 ( .A0N(fu_LSU_wr_mask_x[18]), .A1N(n2247), .B0(n1276), .Y(
        n1012) );
  OAI2BB1X1 U2043 ( .A0N(fu_LSU_wr_mask_x[13]), .A1N(n2248), .B0(n1272), .Y(
        n1008) );
  OAI2BB1X1 U2044 ( .A0N(fu_LSU_wr_mask_x[19]), .A1N(n2247), .B0(n1276), .Y(
        n1015) );
  OAI2BB1X1 U2045 ( .A0N(fu_LSU_wr_mask_x[12]), .A1N(n2248), .B0(n1272), .Y(
        n1003) );
  OAI2BB1X1 U2046 ( .A0N(fu_LSU_wr_mask_x[20]), .A1N(n2248), .B0(n1276), .Y(
        n1011) );
  OAI2BB1X1 U2047 ( .A0N(fu_LSU_wr_mask_x[11]), .A1N(n2248), .B0(n1272), .Y(
        n1007) );
  OAI2BB1X1 U2048 ( .A0N(fu_LSU_wr_mask_x[21]), .A1N(n2247), .B0(n1276), .Y(
        n1016) );
  OAI2BB1X1 U2049 ( .A0N(fu_LSU_wr_mask_x[10]), .A1N(n2248), .B0(n1272), .Y(
        n1004) );
  OAI2BB1X1 U2050 ( .A0N(fu_LSU_wr_mask_x[22]), .A1N(n2248), .B0(n1276), .Y(
        n1010) );
  OAI2BB1X1 U2051 ( .A0N(fu_LSU_wr_mask_x[9]), .A1N(n2248), .B0(n1272), .Y(
        n1006) );
  OAI2BB1X1 U2052 ( .A0N(fu_LSU_wr_mask_x[23]), .A1N(n2247), .B0(n1276), .Y(
        n1017) );
  OAI2BB1X1 U2053 ( .A0N(fu_LSU_wr_mask_x[8]), .A1N(n2248), .B0(n1272), .Y(
        n1005) );
  INVX6 U2054 ( .A(rf_RF_t1data_wire[16]), .Y(n241) );
  CLKNAND2X8 U2055 ( .A(n242), .B(n243), .Y(rf_RF_t1data_wire[16]) );
  INVX6 U2056 ( .A(rf_RF_t1data_wire[17]), .Y(n221) );
  CLKNAND2X8 U2057 ( .A(n222), .B(n223), .Y(rf_RF_t1data_wire[17]) );
  INVX6 U2058 ( .A(rf_RF_t1data_wire[18]), .Y(n208) );
  CLKNAND2X8 U2059 ( .A(n209), .B(n210), .Y(rf_RF_t1data_wire[18]) );
  NAND2X6 U2060 ( .A(n448), .B(n446), .Y(n420) );
  NAND2X2 U2061 ( .A(n2098), .B(n521), .Y(n19) );
  OAI221X2 U2062 ( .A0(n1767), .A1(n2153), .B0(n2059), .B1(
        fu_ALU_fu_arch_sub_200_B_14_), .C0(n2058), .Y(n2060) );
  CLKXOR2X2 U2063 ( .A(n2153), .B(n2154), .Y(n1928) );
  NAND2X5 U2064 ( .A(n206), .B(n1788), .Y(n142) );
  INVX5 U2065 ( .A(n103), .Y(n29) );
  OAI22X4 U2066 ( .A0(n1960), .A1(fu_ALU_o1reg[6]), .B0(n1766), .B1(n2166), 
        .Y(n1966) );
  INVX5 U2067 ( .A(fu_LSU_status_addr_reg_1__2_), .Y(n459) );
  NOR4X4 U2068 ( .A(inst_fetch_reset_cntr_31_), .B(inst_fetch_reset_cntr_30_), 
        .C(inst_fetch_reset_cntr_2_), .D(inst_fetch_reset_cntr_29_), .Y(n614)
         );
  OAI21BX4 U2069 ( .A0(n2271), .A1(n2270), .B0N(inst_fetch_reset_cntr_31_), 
        .Y(inst_fetch_N79) );
  INVX4 U2070 ( .A(rf_RF_t1opcode_wire[0]), .Y(n546) );
  NOR4X4 U2071 ( .A(rf_RF_t1opcode_wire[1]), .B(rf_RF_t1opcode_wire[0]), .C(
        n548), .D(n545), .Y(n47) );
  NOR4X4 U2072 ( .A(rf_RF_t1opcode_wire[2]), .B(rf_RF_t1opcode_wire[0]), .C(
        rf_RF_t1opcode_wire[1]), .D(n545), .Y(n43) );
  NOR4X4 U2073 ( .A(rf_RF_t1opcode_wire[2]), .B(rf_RF_t1opcode_wire[0]), .C(
        n547), .D(n545), .Y(n45) );
  NOR4X4 U2074 ( .A(inst_fetch_reset_cntr_8_), .B(inst_fetch_reset_cntr_7_), 
        .C(inst_fetch_reset_cntr_6_), .D(inst_fetch_reset_cntr_5_), .Y(n2265)
         );
  NOR4X4 U2075 ( .A(inst_fetch_reset_cntr_6_), .B(inst_fetch_reset_cntr_5_), 
        .C(inst_fetch_reset_cntr_4_), .D(inst_fetch_reset_cntr_3_), .Y(n616)
         );
  NOR4X4 U2076 ( .A(inst_fetch_reset_cntr_4_), .B(inst_fetch_reset_cntr_3_), 
        .C(inst_fetch_reset_cntr_30_), .D(inst_fetch_reset_cntr_2_), .Y(n2262)
         );
  NOR4X4 U2077 ( .A(inst_fetch_reset_cntr_21_), .B(inst_fetch_reset_cntr_20_), 
        .C(inst_fetch_reset_cntr_1_), .D(inst_fetch_reset_cntr_19_), .Y(n2269)
         );
  NOR4X4 U2078 ( .A(inst_fetch_reset_cntr_18_), .B(inst_fetch_reset_cntr_17_), 
        .C(inst_fetch_reset_cntr_16_), .D(inst_fetch_reset_cntr_15_), .Y(n2266) );
  NOR4X4 U2079 ( .A(inst_fetch_reset_cntr_29_), .B(inst_fetch_reset_cntr_28_), 
        .C(inst_fetch_reset_cntr_27_), .D(inst_fetch_reset_cntr_26_), .Y(n2263) );
  NOR4X4 U2080 ( .A(inst_fetch_reset_cntr_14_), .B(inst_fetch_reset_cntr_13_), 
        .C(inst_fetch_reset_cntr_12_), .D(inst_fetch_reset_cntr_11_), .Y(n2267) );
  NOR4BX4 U2081 ( .AN(inst_fetch_reset_cntr_0_), .B(inst_fetch_reset_cntr_11_), 
        .C(inst_fetch_reset_cntr_10_), .D(inst_fetch_N79), .Y(n625) );
  NOR3X2 U2082 ( .A(inst_fetch_reset_cntr_10_), .B(inst_fetch_reset_cntr_9_), 
        .C(inst_fetch_reset_cntr_0_), .Y(n2264) );
  NOR4X4 U2083 ( .A(inst_fetch_reset_cntr_13_), .B(inst_fetch_reset_cntr_12_), 
        .C(n618), .D(n619), .Y(n615) );
  NOR4X4 U2084 ( .A(inst_fetch_reset_cntr_25_), .B(inst_fetch_reset_cntr_24_), 
        .C(inst_fetch_reset_cntr_23_), .D(inst_fetch_reset_cntr_22_), .Y(n2268) );
  CLKXOR2X2 U2085 ( .A(fu_ALU_o1reg[6]), .B(n2169), .Y(n1917) );
  NOR4X4 U2086 ( .A(n2182), .B(n239), .C(n132), .D(n2249), .Y(n28) );
  OAI2B11X2 U2087 ( .A1N(fu_ALU_fu_arch_sub_200_B_8_), .A0(n2165), .B0(n1975), 
        .C0(n1982), .Y(n1967) );
  OAI2B11X2 U2088 ( .A1N(fu_ALU_o1reg[8]), .A0(n2165), .B0(n2049), .C0(n2056), 
        .Y(n2041) );
  CLKXOR2X2 U2089 ( .A(fu_ALU_fu_arch_sub_200_B_8_), .B(n2165), .Y(n1930) );
  AOI21X6 U2090 ( .A0(n2197), .A1(fu_ALU_fu_arch_sub_200_B_8_), .B0(
        fu_ALU_fu_arch_n755), .Y(fu_ALU_fu_arch_n157) );
  INVX10 U2091 ( .A(n2164), .Y(fu_ALU_fu_arch_sub_200_B_8_) );
  AOI22X4 U2092 ( .A0(n1775), .A1(fu_ALU_fu_arch_n441), .B0(
        fu_ALU_fu_arch_n249), .B1(n1849), .Y(fu_ALU_fu_arch_n204) );
  BUFX10 U2093 ( .A(n475), .Y(n2118) );
  ADDHX4 U2094 ( .A(inst_fetch_pc_reg_7_), .B(inst_fetch_add_136_carry_7_), 
        .CO(inst_fetch_add_136_carry_8_), .S(inst_fetch_increased_pc_7_) );
  ADDHX4 U2095 ( .A(inst_fetch_pc_reg_8_), .B(inst_fetch_add_136_carry_8_), 
        .CO(inst_fetch_add_136_carry_9_), .S(inst_fetch_increased_pc_8_) );
  ADDHX4 U2096 ( .A(inst_fetch_pc_reg_6_), .B(inst_fetch_add_136_carry_6_), 
        .CO(inst_fetch_add_136_carry_7_), .S(inst_fetch_increased_pc_6_) );
  ADDHX4 U2097 ( .A(inst_fetch_pc_reg_9_), .B(inst_fetch_add_136_carry_9_), 
        .CO(inst_fetch_add_136_carry_10_), .S(inst_fetch_increased_pc_9_) );
  ADDHX4 U2098 ( .A(inst_fetch_pc_reg_5_), .B(inst_fetch_add_136_carry_5_), 
        .CO(inst_fetch_add_136_carry_6_), .S(inst_fetch_increased_pc_5_) );
  ADDHX4 U2099 ( .A(inst_fetch_pc_reg_10_), .B(inst_fetch_add_136_carry_10_), 
        .CO(inst_fetch_add_136_carry_11_), .S(inst_fetch_increased_pc_10_) );
  ADDHX4 U2100 ( .A(inst_fetch_pc_reg_4_), .B(inst_fetch_add_136_carry_4_), 
        .CO(inst_fetch_add_136_carry_5_), .S(inst_fetch_increased_pc_4_) );
  ADDHX4 U2101 ( .A(inst_fetch_pc_reg_11_), .B(inst_fetch_add_136_carry_11_), 
        .CO(inst_fetch_add_136_carry_12_), .S(inst_fetch_increased_pc_11_) );
  ADDHX4 U2102 ( .A(inst_fetch_pc_reg_3_), .B(inst_fetch_add_136_carry_3_), 
        .CO(inst_fetch_add_136_carry_4_), .S(inst_fetch_increased_pc_3_) );
  ADDHX4 U2103 ( .A(inst_fetch_pc_reg_12_), .B(inst_fetch_add_136_carry_12_), 
        .CO(inst_fetch_add_136_carry_13_), .S(inst_fetch_increased_pc_12_) );
  ADDHX4 U2104 ( .A(inst_fetch_pc_reg_2_), .B(inst_fetch_add_136_carry_2_), 
        .CO(inst_fetch_add_136_carry_3_), .S(inst_fetch_increased_pc_2_) );
  ADDHX4 U2105 ( .A(inst_fetch_pc_reg_13_), .B(inst_fetch_add_136_carry_13_), 
        .CO(inst_fetch_add_136_carry_14_), .S(inst_fetch_increased_pc_13_) );
  ADDHX4 U2106 ( .A(inst_fetch_pc_reg_1_), .B(inst_fetch_pc_reg_0_), .CO(
        inst_fetch_add_136_carry_2_), .S(inst_fetch_increased_pc_1_) );
  BUFX12 U2107 ( .A(n2221), .Y(n2222) );
  BUFX16 U2108 ( .A(n52), .Y(n2221) );
  CLKXOR2X2 U2109 ( .A(n2157), .B(n2158), .Y(n1929) );
  CLKXOR2X2 U2110 ( .A(n2136), .B(n2137), .Y(n1912) );
  NAND3X4 U2111 ( .A(n543), .B(inst_decoder_instructionword_wire[4]), .C(n551), 
        .Y(n538) );
  NAND2BX4 U2112 ( .AN(inst_decoder_instructionword_wire[4]), .B(n566), .Y(
        n552) );
  OAI211X2 U2113 ( .A0(inst_decoder_instructionword_wire[40]), .A1(n557), .B0(
        n595), .C0(n596), .Y(n594) );
  CLKBUFX6 U2114 ( .A(n463), .Y(n1863) );
  INVX6 U2115 ( .A(n320), .Y(n252) );
  BUFX12 U2116 ( .A(n1777), .Y(n2214) );
  INVX4 U2117 ( .A(fu_ALU_o1reg[4]), .Y(n2171) );
  BUFX10 U2118 ( .A(n2094), .Y(n2203) );
  OR2X2 U2119 ( .A(n2174), .B(fu_ALU_fu_arch_n335), .Y(n2094) );
  BUFX10 U2120 ( .A(fu_ALU_fu_arch_n394), .Y(n2101) );
  AOI2B1X4 U2121 ( .A1N(n2179), .A0(fu_ALU_fu_arch_sub_200_B_14_), .B0(n2046), 
        .Y(n2062) );
  CLKXOR2X2 U2122 ( .A(fu_ALU_fu_arch_sub_200_B_14_), .B(n2179), .Y(n1921) );
  XNOR2X2 U2123 ( .A(n2180), .B(fu_ALU_o1reg[31]), .Y(n1914) );
  CLKXOR2X2 U2124 ( .A(fu_ALU_o1reg[20]), .B(n2145), .Y(n1905) );
  AOI2B1X4 U2125 ( .A1N(n2126), .A0(fu_ALU_fu_arch_sub_200_B_30_), .B0(n1943), 
        .Y(n1954) );
  XNOR2X2 U2126 ( .A(fu_ALU_fu_arch_sub_200_B_30_), .B(n2126), .Y(n1915) );
  NOR3X4 U2127 ( .A(n2212), .B(fu_LSU_status_addr_reg_1__4_), .C(
        fu_LSU_status_addr_reg_1__3_), .Y(n475) );
  INVX5 U2128 ( .A(inst_decoder_N230), .Y(n537) );
  INVX4 U2129 ( .A(fu_LSU_t1opcode_wire[1]), .Y(n239) );
  OAI21X6 U2130 ( .A0(n2183), .A1(fu_LSU_t1opcode_wire[1]), .B0(
        fu_LSU_t1opcode_wire[2]), .Y(n417) );
  NOR2X3 U2131 ( .A(n2183), .B(fu_LSU_t1opcode_wire[1]), .Y(n526) );
  OAI31X4 U2132 ( .A0(n1806), .A1(n2212), .A2(n493), .B0(n462), .Y(n472) );
  BUFX12 U2133 ( .A(n267), .Y(n2116) );
  BUFX12 U2134 ( .A(n2250), .Y(n2251) );
  INVX4 U2135 ( .A(inst_decoder_instructionword_wire[35]), .Y(n578) );
  INVX4 U2136 ( .A(fu_ALU_opc1reg[2]), .Y(fu_ALU_fu_arch_n760) );
  NOR4X4 U2137 ( .A(fu_ALU_opc1reg[0]), .B(fu_ALU_opc1reg[2]), .C(
        fu_ALU_opc1reg[3]), .D(fu_ALU_opc1reg[1]), .Y(fu_ALU_fu_arch_n130) );
  NOR4X4 U2138 ( .A(fu_ALU_opc1reg[2]), .B(fu_ALU_opc1reg[3]), .C(
        fu_ALU_fu_arch_n752), .D(fu_ALU_fu_arch_n744), .Y(fu_ALU_fu_arch_n747)
         );
  INVX4 U2139 ( .A(fu_ALU_opc1reg[1]), .Y(fu_ALU_fu_arch_n744) );
  NOR3X4 U2140 ( .A(fu_ALU_opc1reg[1]), .B(fu_ALU_fu_arch_n746), .C(
        fu_ALU_fu_arch_n745), .Y(fu_ALU_fu_arch_n129) );
  CLKINVX24 U2141 ( .A(n2098), .Y(n2253) );
  BUFX12 U2142 ( .A(n2248), .Y(n2247) );
  CLKBUFX40 U2143 ( .A(n32), .Y(n2248) );
  INVX2 U2144 ( .A(fu_ALU_o1reg[24]), .Y(fu_ALU_fu_arch_sub_200_B_not_24_) );
  INVX4 U2145 ( .A(fu_ALU_o1reg[11]), .Y(n2159) );
  INVX4 U2146 ( .A(rstx), .Y(n2261) );
  INVX4 U2147 ( .A(rstx), .Y(n2260) );
  NAND2X4 U2148 ( .A(rf_BOOL_t1opcode_wire_0_), .B(rf_BOOL_t1load_wire), .Y(
        n605) );
  INVX4 U2149 ( .A(fu_ALU_t1reg[5]), .Y(n2039) );
  INVX4 U2150 ( .A(fu_ALU_fu_arch_n278), .Y(fu_ALU_fu_arch_n308) );
  INVX4 U2151 ( .A(fu_LSU_t1opcode_wire[2]), .Y(n527) );
  INVX4 U2152 ( .A(inst_decoder_instructionword_wire[37]), .Y(n579) );
  CLKBUFX32 U2153 ( .A(ic_socket_LIFTING_o1_bus_cntrl_wire_0_), .Y(n2256) );
  AOI221X2 U2154 ( .A0(n2186), .A1(ic_socket_gcu_o1_data0_wire[1]), .B0(n2257), 
        .B1(ic_socket_ALU_o1_data0_wire[1]), .C0(n632), .Y(n627) );
  CLKBUFX32 U2155 ( .A(ic_socket_ALU_o1_bus_cntrl_wire_0_), .Y(n2257) );
  NOR2X3 U2156 ( .A(n2150), .B(n2195), .Y(fu_ALU_fu_arch_n598) );
  OAI211X2 U2157 ( .A0(fu_ALU_fu_arch_n462), .A1(fu_ALU_fu_arch_n463), .B0(
        fu_ALU_fu_arch_n464), .C0(fu_ALU_fu_arch_n465), .Y(
        ic_socket_ALU_o1_data0_wire[23]) );
  OAI211X2 U2158 ( .A0(fu_ALU_fu_arch_n483), .A1(fu_ALU_fu_arch_n463), .B0(
        fu_ALU_fu_arch_n484), .C0(fu_ALU_fu_arch_n485), .Y(
        ic_socket_ALU_o1_data0_wire[22]) );
  INVX4 U2159 ( .A(n2100), .Y(fu_ALU_fu_arch_n463) );
  OAI211X2 U2160 ( .A0(n1776), .A1(fu_ALU_fu_arch_n621), .B0(
        fu_ALU_fu_arch_n623), .C0(fu_ALU_fu_arch_n589), .Y(fu_ALU_fu_arch_n756) );
  CLKXOR2X2 U2161 ( .A(fu_ALU_fu_arch_sub_200_B_5_), .B(fu_ALU_t1reg[5]), .Y(
        n1924) );
  NOR4X4 U2162 ( .A(n1939), .B(n1938), .C(n1937), .D(n1936), .Y(n1940) );
  NOR4X4 U2163 ( .A(n1920), .B(n1919), .C(n1918), .D(n1917), .Y(n1935) );
  NOR4X4 U2164 ( .A(n1927), .B(n1926), .C(n1925), .D(n1924), .Y(n1933) );
  CLKXOR2X2 U2165 ( .A(fu_ALU_fu_arch_sub_200_B_9_), .B(n2163), .Y(n1926) );
  NOR4X4 U2166 ( .A(n1931), .B(n1930), .C(n1929), .D(n1928), .Y(n1932) );
  OAI2B11X2 U2167 ( .A1N(fu_ALU_fu_arch_n229), .A0(fu_ALU_fu_arch_n118), .B0(
        fu_ALU_fu_arch_n230), .C0(fu_ALU_fu_arch_n231), .Y(
        ic_socket_ALU_o1_data0_wire[3]) );
  INVX2 U2168 ( .A(n1879), .Y(n1880) );
  OAI211X2 U2169 ( .A0(n1880), .A1(fu_ALU_fu_arch_n388), .B0(
        fu_ALU_fu_arch_n476), .C0(fu_ALU_fu_arch_n477), .Y(fu_ALU_fu_arch_n470) );
  NAND2X3 U2170 ( .A(n417), .B(n2113), .Y(n501) );
  AOI211X2 U2171 ( .A0(n2028), .A1(n2027), .B0(n2026), .C0(n2025), .Y(n2091)
         );
  NOR4X4 U2172 ( .A(n1923), .B(n1922), .C(fu_ALU_fu_arch_N33), .D(n1921), .Y(
        n1934) );
  NOR4X4 U2173 ( .A(n1913), .B(n1912), .C(n1911), .D(n1910), .Y(n1916) );
  CLKINVX24 U2174 ( .A(n2259), .Y(n2258) );
  CLKNAND2X12 U2175 ( .A(n239), .B(n2117), .Y(n25) );
  BUFX12 U2176 ( .A(n2096), .Y(n2117) );
  NOR2BX4 U2177 ( .AN(n1780), .B(n2135), .Y(n2087) );
  BUFX12 U2178 ( .A(n275), .Y(n2114) );
  NOR2X4 U2179 ( .A(n2109), .B(n1764), .Y(fu_ALU_fu_arch_n310) );
  OAI211X2 U2180 ( .A0(fu_ALU_fu_arch_n607), .A1(n1797), .B0(
        fu_ALU_fu_arch_n609), .C0(fu_ALU_fu_arch_n610), .Y(
        ic_socket_ALU_o1_data0_wire[16]) );
  OAI211X4 U2181 ( .A0(fu_ALU_fu_arch_n499), .A1(n2203), .B0(
        fu_ALU_fu_arch_n727), .C0(fu_ALU_fu_arch_n437), .Y(fu_ALU_fu_arch_n405) );
  AOI2B1X4 U2182 ( .A1N(n2162), .A0(n2161), .B0(n1978), .Y(n1982) );
  AOI2B1X4 U2183 ( .A1N(n2162), .A0(n2161), .B0(n2052), .Y(n2056) );
  NOR2X8 U2184 ( .A(inst_fetch_reset_lock), .B(busy), .Y(n498) );
  AOI222X4 U2185 ( .A0(n1849), .A1(n1775), .B0(n1837), .B1(fu_ALU_fu_arch_n249), .C0(fu_ALU_fu_arch_n441), .C1(n2104), .Y(fu_ALU_fu_arch_n107) );
  CLKNAND2X8 U2186 ( .A(n1883), .B(n1884), .Y(rf_RF_t1data_wire[11]) );
  AOI221X2 U2187 ( .A0(n2186), .A1(ic_socket_gcu_o1_data0_wire[11]), .B0(n2257), .B1(ic_socket_ALU_o1_data0_wire[11]), .C0(n304), .Y(n300) );
  CLKNAND2X8 U2188 ( .A(n1885), .B(n1886), .Y(rf_RF_t1data_wire[14]) );
  AOI221X2 U2189 ( .A0(n2186), .A1(ic_socket_gcu_o1_data0_wire[14]), .B0(n2257), .B1(ic_socket_ALU_o1_data0_wire[14]), .C0(n511), .Y(n507) );
  INVX4 U2190 ( .A(rf_RF_t1opcode_wire[1]), .Y(n547) );
  AOI22X4 U2191 ( .A0(n2176), .A1(fu_ALU_fu_arch_n619), .B0(n1887), .B1(
        fu_ALU_fu_arch_n335), .Y(fu_ALU_fu_arch_n533) );
  CLKBUFX4 U2192 ( .A(fu_ALU_fu_arch_n493), .Y(n1888) );
  AOI222X4 U2193 ( .A0(n1843), .A1(n1775), .B0(n1888), .B1(fu_ALU_fu_arch_n249), .C0(fu_ALU_fu_arch_n334), .C1(n2104), .Y(fu_ALU_fu_arch_n408) );
  OAI211X2 U2194 ( .A0(n1778), .A1(n1776), .B0(fu_ALU_fu_arch_n724), .C0(
        fu_ALU_fu_arch_n327), .Y(fu_ALU_fu_arch_n493) );
  CLKBUFX24 U2195 ( .A(n39), .Y(n2245) );
  AOI22X4 U2196 ( .A0(n1775), .A1(fu_ALU_fu_arch_n434), .B0(
        fu_ALU_fu_arch_n249), .B1(fu_ALU_fu_arch_n435), .Y(fu_ALU_fu_arch_n117) );
  INVX4 U2197 ( .A(n1892), .Y(fu_ALU_fu_arch_n132) );
  INVX2 U2198 ( .A(inst_decoder_instructionword_wire[37]), .Y(n1895) );
  INVX2 U2199 ( .A(inst_decoder_instructionword_wire[36]), .Y(n1896) );
  INVX2 U2200 ( .A(n2183), .Y(n1897) );
  INVX4 U2201 ( .A(fu_LSU_status_addr_reg_1__3_), .Y(n458) );
  CLKXOR2X2 U2202 ( .A(fu_ALU_o1reg[23]), .B(n2139), .Y(n1904) );
  CLKXOR2X2 U2203 ( .A(fu_ALU_o1reg[22]), .B(n2141), .Y(n1903) );
  AOI22X2 U2204 ( .A0(fu_ALU_opc1reg[0]), .A1(fu_ALU_fu_arch_N98), .B0(
        fu_ALU_fu_arch_N97), .B1(fu_ALU_fu_arch_n746), .Y(fu_ALU_fu_arch_n752)
         );
  NAND2X4 U2205 ( .A(fu_ALU_opc1reg[3]), .B(fu_ALU_fu_arch_n760), .Y(
        fu_ALU_fu_arch_n745) );
  OR3X2 U2206 ( .A(fu_ALU_fu_arch_n760), .B(fu_ALU_fu_arch_n744), .C(
        fu_ALU_opc1reg[3]), .Y(fu_ALU_fu_arch_n761) );
  AOI2BB1X4 U2207 ( .A0N(n454), .A1N(n455), .B0(n456), .Y(n452) );
  INVX8 U2208 ( .A(fu_LSU_status_addr_reg_1__1_), .Y(n446) );
  NOR2BX1 U2209 ( .AN(n2180), .B(n2124), .Y(n1943) );
  OAI22X1 U2210 ( .A0(n1944), .A1(fu_ALU_fu_arch_lt_gt_188_A_28_), .B0(n1765), 
        .B1(fu_ALU_fu_arch_sub_200_B_29_), .Y(n1953) );
  AOI2B1X1 U2211 ( .A1N(n1780), .A0(n2135), .B0(n1946), .Y(n1949) );
  OAI2BB1X1 U2212 ( .A0N(n1774), .A1N(n2180), .B0(n2126), .Y(n1950) );
  OAI22X1 U2213 ( .A0(n1955), .A1(n2181), .B0(n1770), .B1(n2177), .Y(n1957) );
  NOR2BX1 U2214 ( .AN(n2153), .B(n2154), .Y(n1972) );
  OAI2BB1X1 U2215 ( .A0N(n1767), .A1N(n2153), .B0(n2179), .Y(n1985) );
  NAND2BX1 U2216 ( .AN(fu_ALU_fu_arch_sub_200_B_9_), .B(n2163), .Y(n1976) );
  AOI21X1 U2217 ( .A0(n1977), .A1(n1976), .B0(n1980), .Y(n1983) );
  AOI2B1X1 U2218 ( .A1N(fu_ALU_fu_arch_sub_200_B_11_), .A0(n2160), .B0(n1979), 
        .Y(n1981) );
  NOR2BX1 U2219 ( .AN(n2151), .B(n2152), .Y(n1994) );
  NOR2BX1 U2220 ( .AN(n2138), .B(n2139), .Y(n1991) );
  NAND2BX2 U2221 ( .AN(n2147), .B(fu_ALU_fu_arch_sub_200_B_19_), .Y(n1999) );
  OAI2BB1X1 U2222 ( .A0N(n1736), .A1N(fu_ALU_fu_arch_sub_200_B_21_), .B0(n2145), .Y(n1996) );
  OAI22X1 U2223 ( .A0(n1996), .A1(n2144), .B0(n1736), .B1(
        fu_ALU_fu_arch_sub_200_B_21_), .Y(n2007) );
  AOI2B1X1 U2224 ( .A1N(fu_ALU_o1reg[17]), .A0(n2150), .B0(n1998), .Y(n2001)
         );
  NOR2BX1 U2225 ( .AN(n2136), .B(n2137), .Y(n2010) );
  OAI2BB1X1 U2226 ( .A0N(n1765), .A1N(fu_ALU_fu_arch_sub_200_B_29_), .B0(n2130), .Y(n1944) );
  NAND2BX2 U2227 ( .AN(n2131), .B(fu_ALU_fu_arch_sub_200_B_27_), .Y(n1947) );
  AOI32X1 U2228 ( .A0(n1763), .A1(n1947), .A2(n2133), .B0(n2131), .B1(n1764), 
        .Y(n1948) );
  OAI2BB1X1 U2229 ( .A0N(n1768), .A1N(n2173), .B0(n2176), .Y(n1959) );
  OAI2BB1X1 U2230 ( .A0N(n1770), .A1N(n2177), .B0(n1779), .Y(n1955) );
  NAND2BX1 U2231 ( .AN(n2176), .B(fu_ALU_fu_arch_sub_200_B_2_), .Y(n1956) );
  OAI2B11X1 U2232 ( .A1N(n2173), .A0(n2174), .B0(n1957), .C0(n1956), .Y(n1958)
         );
  NAND2BX1 U2233 ( .AN(n2172), .B(fu_ALU_fu_arch_sub_200_B_4_), .Y(n1961) );
  OAI2BB1X1 U2234 ( .A0N(n1766), .A1N(n2166), .B0(n2169), .Y(n1960) );
  AOI31X1 U2235 ( .A0(n1963), .A1(n1962), .A2(n1961), .B0(n1966), .Y(n1971) );
  OAI2BB1X1 U2236 ( .A0N(n1965), .A1N(fu_ALU_fu_arch_sub_200_B_5_), .B0(n2172), 
        .Y(n1964) );
  NAND2BX2 U2237 ( .AN(n2163), .B(fu_ALU_fu_arch_sub_200_B_9_), .Y(n1975) );
  AOI221X2 U2238 ( .A0(n1971), .A1(n1970), .B0(n1969), .B1(n1968), .C0(n1967), 
        .Y(n1990) );
  OAI2B11X4 U2239 ( .A1N(fu_ALU_o1reg[13]), .A0(n2156), .B0(n1973), .C0(n1988), 
        .Y(n1980) );
  OAI2BB1X1 U2240 ( .A0N(n1740), .A1N(fu_ALU_o1reg[13]), .B0(n2158), .Y(n1974)
         );
  NAND3BX1 U2241 ( .AN(fu_ALU_fu_arch_sub_200_B_8_), .B(n1975), .C(n2165), .Y(
        n1977) );
  AOI221X2 U2242 ( .A0(n1990), .A1(n1989), .B0(n1988), .B1(n1987), .C0(n1986), 
        .Y(n1995) );
  NAND2BX1 U2243 ( .AN(n2145), .B(n2144), .Y(n1992) );
  AOI32X1 U2244 ( .A0(n1771), .A1(n1999), .A2(n2149), .B0(n2147), .B1(n2146), 
        .Y(n2000) );
  OAI2BB1X1 U2245 ( .A0N(n1737), .A1N(n2138), .B0(n2141), .Y(n2004) );
  AOI32X2 U2246 ( .A0(n1787), .A1(n2015), .A2(n2014), .B0(n2013), .B1(n1787), 
        .Y(fu_ALU_fu_arch_N98) );
  OR4X2 U2247 ( .A(n1997), .B(n1995), .C(n1994), .D(n1993), .Y(n2015) );
  AOI2B1X4 U2248 ( .A1N(n2179), .A0(fu_ALU_fu_arch_sub_200_B_14_), .B0(n1972), 
        .Y(n1988) );
  OAI221X2 U2249 ( .A0(n1767), .A1(n2153), .B0(n1985), .B1(
        fu_ALU_fu_arch_sub_200_B_14_), .C0(n1984), .Y(n1986) );
  AOI2B1X4 U2250 ( .A1N(n2141), .A0(fu_ALU_o1reg[22]), .B0(n1991), .Y(n2008)
         );
  NOR2BX4 U2251 ( .AN(n1780), .B(n2135), .Y(n2012) );
  NAND2BX2 U2252 ( .AN(n2158), .B(n2157), .Y(n1973) );
  INVX2 U2253 ( .A(n1980), .Y(n1989) );
  NOR2BX1 U2254 ( .AN(n2124), .B(n2180), .Y(n2017) );
  OAI22X1 U2255 ( .A0(n2018), .A1(fu_ALU_fu_arch_lt_gt_188_A_28_), .B0(n1765), 
        .B1(fu_ALU_fu_arch_sub_200_B_29_), .Y(n2027) );
  AOI2B1X1 U2256 ( .A1N(n1780), .A0(n2135), .B0(n2020), .Y(n2023) );
  OAI2BB1X1 U2257 ( .A0N(n1739), .A1N(n2124), .B0(n2126), .Y(n2024) );
  OAI22X1 U2258 ( .A0(n2024), .A1(fu_ALU_fu_arch_sub_200_B_30_), .B0(n1739), 
        .B1(n2124), .Y(n2025) );
  OAI22X1 U2259 ( .A0(n2029), .A1(n2181), .B0(n1770), .B1(n2177), .Y(n2031) );
  NAND2BX1 U2260 ( .AN(n2158), .B(n2157), .Y(n2047) );
  NOR2BX1 U2261 ( .AN(n2153), .B(n2154), .Y(n2046) );
  OAI22X1 U2262 ( .A0(n2048), .A1(n2157), .B0(n1740), .B1(fu_ALU_o1reg[13]), 
        .Y(n2061) );
  OAI2BB1X1 U2263 ( .A0N(n1767), .A1N(n2153), .B0(n2179), .Y(n2059) );
  NAND2BX1 U2264 ( .AN(fu_ALU_fu_arch_sub_200_B_9_), .B(n2163), .Y(n2050) );
  AOI21X1 U2265 ( .A0(n2051), .A1(n2050), .B0(n1783), .Y(n2057) );
  AOI2B1X1 U2266 ( .A1N(fu_ALU_fu_arch_sub_200_B_11_), .A0(n2160), .B0(n2053), 
        .Y(n2055) );
  NOR2BX1 U2267 ( .AN(n2151), .B(n2152), .Y(n2068) );
  NOR2BX1 U2268 ( .AN(n2138), .B(n2139), .Y(n2065) );
  OAI2BB1X1 U2269 ( .A0N(n1736), .A1N(fu_ALU_fu_arch_sub_200_B_21_), .B0(n2145), .Y(n2070) );
  OAI22X1 U2270 ( .A0(n2070), .A1(n2144), .B0(n1736), .B1(
        fu_ALU_fu_arch_sub_200_B_21_), .Y(n2082) );
  AOI2B1X1 U2271 ( .A1N(fu_ALU_o1reg[17]), .A0(n2150), .B0(n2072), .Y(n2076)
         );
  OAI22X1 U2272 ( .A0(n2079), .A1(fu_ALU_fu_arch_sub_200_B_22_), .B0(n1737), 
        .B1(n2138), .Y(n2080) );
  NOR2BX1 U2273 ( .AN(n2136), .B(n2137), .Y(n2085) );
  OAI2BB1X1 U2274 ( .A0N(n1765), .A1N(fu_ALU_fu_arch_sub_200_B_29_), .B0(n2130), .Y(n2018) );
  NAND2BX2 U2275 ( .AN(n2131), .B(fu_ALU_fu_arch_sub_200_B_27_), .Y(n2021) );
  AOI32X1 U2276 ( .A0(n1763), .A1(n2021), .A2(n2133), .B0(n2131), .B1(n1764), 
        .Y(n2022) );
  OAI2BB1X1 U2277 ( .A0N(n1768), .A1N(n2173), .B0(n2176), .Y(n2033) );
  OAI2BB1X1 U2278 ( .A0N(n1770), .A1N(n2177), .B0(n1779), .Y(n2029) );
  NAND2BX1 U2279 ( .AN(n2176), .B(fu_ALU_fu_arch_sub_200_B_2_), .Y(n2030) );
  OAI2B11X1 U2280 ( .A1N(n2173), .A0(n2174), .B0(n2031), .C0(n2030), .Y(n2032)
         );
  NAND2BX1 U2281 ( .AN(n2172), .B(fu_ALU_o1reg[4]), .Y(n2035) );
  OAI2BB1X1 U2282 ( .A0N(n1766), .A1N(n2166), .B0(n2169), .Y(n2034) );
  AOI31X1 U2283 ( .A0(n2037), .A1(n2036), .A2(n2035), .B0(n2040), .Y(n2045) );
  OAI2BB1X1 U2284 ( .A0N(n2039), .A1N(fu_ALU_fu_arch_sub_200_B_5_), .B0(n2172), 
        .Y(n2038) );
  NAND2BX2 U2285 ( .AN(n2163), .B(fu_ALU_fu_arch_sub_200_B_9_), .Y(n2049) );
  AOI221X2 U2286 ( .A0(n2045), .A1(n2044), .B0(n2043), .B1(n2042), .C0(n2041), 
        .Y(n2064) );
  OAI2BB1X1 U2287 ( .A0N(n1740), .A1N(fu_ALU_o1reg[13]), .B0(n2158), .Y(n2048)
         );
  NAND3BX1 U2288 ( .AN(fu_ALU_o1reg[8]), .B(n2049), .C(n2165), .Y(n2051) );
  AOI221X2 U2289 ( .A0(n2064), .A1(n2063), .B0(n2062), .B1(n2061), .C0(n2060), 
        .Y(n2069) );
  NAND2BX2 U2290 ( .AN(n2147), .B(fu_ALU_o1reg[19]), .Y(n2074) );
  CLKINVX1 U2291 ( .A(fu_ALU_o1reg[19]), .Y(n2073) );
  AOI32X1 U2292 ( .A0(n1771), .A1(n2074), .A2(n2149), .B0(n2147), .B1(n2073), 
        .Y(n2075) );
  OAI2BB1X1 U2293 ( .A0N(n1737), .A1N(n2138), .B0(n2141), .Y(n2079) );
  NOR3BX2 U2294 ( .AN(n2162), .B(n2052), .C(n2161), .Y(n2053) );
  AOI2B1X4 U2295 ( .A1N(n2126), .A0(fu_ALU_fu_arch_sub_200_B_30_), .B0(n2017), 
        .Y(n2028) );
  OR4X2 U2296 ( .A(n2071), .B(n2069), .C(n2068), .D(n2067), .Y(n2090) );
  AOI2B1X4 U2297 ( .A1N(n2141), .A0(fu_ALU_fu_arch_sub_200_B_22_), .B0(n2065), 
        .Y(n2083) );
  NAND2BX2 U2298 ( .AN(n2145), .B(n2144), .Y(n2066) );
  CLKXOR2X2 U2299 ( .A(inst_fetch_add_136_carry_14_), .B(inst_fetch_pc_reg_14_), .Y(inst_fetch_increased_pc_14_) );
  BUFX8 U2300 ( .A(fu_ALU_fu_arch_n352), .Y(n2102) );
  AND4X4 U2301 ( .A(n627), .B(n628), .C(n629), .D(n630), .Y(n2096) );
  CLKBUFX4 U2302 ( .A(n2193), .Y(n2194) );
  INVX8 U2303 ( .A(n2104), .Y(fu_ALU_fu_arch_n468) );
  INVX10 U2304 ( .A(n1754), .Y(fu_ALU_fu_arch_sub_200_B_5_) );
  CLKINVX40 U2305 ( .A(n2092), .Y(n2190) );
  BUFX12 U2306 ( .A(n2191), .Y(n2192) );
  CLKINVX24 U2307 ( .A(n2207), .Y(n2206) );
  CLKNAND2X8 U2308 ( .A(n2172), .B(fu_ALU_fu_arch_n274), .Y(
        fu_ALU_fu_arch_n212) );
  CLKBUFX24 U2309 ( .A(fu_ALU_fu_arch_n284), .Y(n2202) );
  INVX18 U2310 ( .A(n1762), .Y(n2195) );
  INVX4 U2311 ( .A(fu_ALU_o1reg[28]), .Y(n2129) );
  CLKNAND2X8 U2312 ( .A(fu_ALU_fu_arch_n274), .B(fu_ALU_fu_arch_n220), .Y(
        fu_ALU_fu_arch_n292) );
  BUFX10 U2313 ( .A(fu_ALU_fu_arch_n379), .Y(n2106) );
  CLKBUFX6 U2314 ( .A(n57), .Y(n2218) );
  NOR3X2 U2315 ( .A(n584), .B(n1748), .C(n582), .Y(n57) );
  CLKINVX32 U2316 ( .A(n2098), .Y(n2252) );
  BUFX10 U2317 ( .A(n53), .Y(n2220) );
  CLKBUFX24 U2318 ( .A(n2095), .Y(n2201) );
  CLKBUFX16 U2319 ( .A(n53), .Y(n2219) );
  OAI22X1 fu_LIFTING_U613 ( .A0(fu_LIFTING_n46), .A1(fu_LIFTING_n1), .B0(
        fu_LIFTING_n45), .B1(fu_LIFTING_n237), .Y(fu_LIFTING_n273) );
  OAI22X1 fu_LIFTING_U612 ( .A0(fu_LIFTING_n47), .A1(fu_LIFTING_n1), .B0(
        fu_LIFTING_n48), .B1(fu_LIFTING_n237), .Y(fu_LIFTING_n276) );
  OAI22X1 fu_LIFTING_U611 ( .A0(fu_LIFTING_n63), .A1(fu_LIFTING_n1), .B0(
        fu_LIFTING_n62), .B1(fu_LIFTING_n237), .Y(fu_LIFTING_n309) );
  OAI22X1 fu_LIFTING_U610 ( .A0(fu_LIFTING_n68), .A1(fu_LIFTING_n1), .B0(
        fu_LIFTING_n69), .B1(fu_LIFTING_n237), .Y(fu_LIFTING_n324) );
  OAI22X1 fu_LIFTING_U609 ( .A0(fu_LIFTING_n73), .A1(fu_LIFTING_n2), .B0(
        fu_LIFTING_n339), .B1(fu_LIFTING_n237), .Y(fu_LIFTING_n340) );
  OAI22X1 fu_LIFTING_U608 ( .A0(fu_LIFTING_n354), .A1(fu_LIFTING_n2), .B0(
        fu_LIFTING_n39), .B1(fu_LIFTING_n237), .Y(fu_LIFTING_n351) );
  OAI21X1 fu_LIFTING_U607 ( .A0(fu_LIFTING_n36), .A1(fu_LIFTING_n234), .B0(
        fu_LIFTING_N72), .Y(fu_LIFTING_n260) );
  CLKMX2X12 fu_LIFTING_U606 ( .A(fu_LIFTING_reg_x1_24_), .B(
        rf_RF_t1data_wire[24]), .S0(fu_LIFTING_n249), .Y(fu_LIFTING_N79) );
  CLKMX2X12 fu_LIFTING_U605 ( .A(fu_LIFTING_reg_x1_18_), .B(
        rf_RF_t1data_wire[18]), .S0(fu_LIFTING_n42), .Y(fu_LIFTING_N85) );
  CLKMX2X12 fu_LIFTING_U604 ( .A(fu_LIFTING_reg_x1_15_), .B(
        rf_RF_t1data_wire[15]), .S0(fu_LIFTING_n42), .Y(fu_LIFTING_N88) );
  CLKMX2X12 fu_LIFTING_U603 ( .A(fu_LIFTING_reg_x1_14_), .B(
        rf_RF_t1data_wire[14]), .S0(fu_LIFTING_n42), .Y(fu_LIFTING_N89) );
  CLKMX2X12 fu_LIFTING_U602 ( .A(fu_LIFTING_reg_x1_13_), .B(n1823), .S0(
        fu_LIFTING_n42), .Y(fu_LIFTING_N90) );
  CLKMX2X12 fu_LIFTING_U601 ( .A(fu_LIFTING_reg_x1_10_), .B(n1816), .S0(
        fu_LIFTING_n42), .Y(fu_LIFTING_N93) );
  CLKMX2X12 fu_LIFTING_U600 ( .A(fu_LIFTING_reg_x1_4_), .B(n1825), .S0(
        fu_LIFTING_n42), .Y(fu_LIFTING_N99) );
  CLKMX2X12 fu_LIFTING_U599 ( .A(fu_LIFTING_reg_x2_24_), .B(
        rf_RF_t1data_wire[24]), .S0(fu_LIFTING_n248), .Y(fu_LIFTING_N679) );
  CLKMX2X12 fu_LIFTING_U598 ( .A(fu_LIFTING_reg_x2_18_), .B(
        rf_RF_t1data_wire[18]), .S0(fu_LIFTING_n248), .Y(fu_LIFTING_N685) );
  CLKMX2X12 fu_LIFTING_U597 ( .A(fu_LIFTING_reg_x2_15_), .B(
        rf_RF_t1data_wire[15]), .S0(fu_LIFTING_n248), .Y(fu_LIFTING_N688) );
  CLKMX2X12 fu_LIFTING_U596 ( .A(fu_LIFTING_reg_x2_13_), .B(n1823), .S0(
        fu_LIFTING_n248), .Y(fu_LIFTING_N690) );
  CLKMX2X12 fu_LIFTING_U595 ( .A(fu_LIFTING_reg_x2_10_), .B(n1816), .S0(
        fu_LIFTING_n248), .Y(fu_LIFTING_N693) );
  CLKMX2X12 fu_LIFTING_U594 ( .A(fu_LIFTING_reg_x2_6_), .B(n1818), .S0(
        fu_LIFTING_n248), .Y(fu_LIFTING_N697) );
  CLKMX2X12 fu_LIFTING_U593 ( .A(fu_LIFTING_reg_x2_5_), .B(
        rf_RF_t1data_wire[5]), .S0(fu_LIFTING_n248), .Y(fu_LIFTING_N698) );
  CLKMX2X12 fu_LIFTING_U592 ( .A(fu_LIFTING_reg_x2_3_), .B(
        rf_RF_t1data_wire[3]), .S0(fu_LIFTING_n248), .Y(fu_LIFTING_N700) );
  CLKMX2X12 fu_LIFTING_U591 ( .A(fu_LIFTING_reg_x2_1_), .B(n2110), .S0(
        fu_LIFTING_n248), .Y(fu_LIFTING_N702) );
  AOI222X4 fu_LIFTING_U590 ( .A0(fu_LIFTING_N671), .A1(fu_LIFTING_n240), .B0(
        fu_LIFTING_n234), .B1(fu_LIFTING_N311), .C0(fu_LIFTING_n238), .C1(
        fu_LIFTING_N191), .Y(fu_LIFTING_n362) );
  AOI222X4 fu_LIFTING_U589 ( .A0(fu_LIFTING_N71), .A1(fu_LIFTING_n36), .B0(
        fu_LIFTING_n83), .B1(fu_LIFTING_N431), .C0(fu_LIFTING_n37), .C1(
        fu_LIFTING_N551), .Y(fu_LIFTING_n361) );
  AOI21X1 fu_LIFTING_U588 ( .A0(fu_LIFTING_n241), .A1(fu_LIFTING_n239), .B0(
        fu_LIFTING_n266), .Y(fu_LIFTING_n263) );
  AOI21X1 fu_LIFTING_U587 ( .A0(fu_LIFTING_n37), .A1(fu_LIFTING_N73), .B0(
        fu_LIFTING_n263), .Y(fu_LIFTING_n265) );
  OAI21X1 fu_LIFTING_U586 ( .A0(fu_LIFTING_n36), .A1(fu_LIFTING_n234), .B0(
        fu_LIFTING_N73), .Y(fu_LIFTING_n264) );
  AOI21X1 fu_LIFTING_U585 ( .A0(fu_LIFTING_n241), .A1(fu_LIFTING_n239), .B0(
        fu_LIFTING_n43), .Y(fu_LIFTING_n267) );
  OAI21X1 fu_LIFTING_U584 ( .A0(fu_LIFTING_n36), .A1(fu_LIFTING_n234), .B0(
        fu_LIFTING_N74), .Y(fu_LIFTING_n268) );
  AOI21X1 fu_LIFTING_U583 ( .A0(fu_LIFTING_n241), .A1(fu_LIFTING_n239), .B0(
        fu_LIFTING_n44), .Y(fu_LIFTING_n270) );
  AOI21X1 fu_LIFTING_U582 ( .A0(fu_LIFTING_n37), .A1(fu_LIFTING_N75), .B0(
        fu_LIFTING_n270), .Y(fu_LIFTING_n272) );
  OAI21X1 fu_LIFTING_U581 ( .A0(fu_LIFTING_n36), .A1(fu_LIFTING_n234), .B0(
        fu_LIFTING_N75), .Y(fu_LIFTING_n271) );
  AOI21X1 fu_LIFTING_U580 ( .A0(fu_LIFTING_n36), .A1(fu_LIFTING_N76), .B0(
        fu_LIFTING_n273), .Y(fu_LIFTING_n275) );
  AOI21X1 fu_LIFTING_U579 ( .A0(fu_LIFTING_n36), .A1(fu_LIFTING_N77), .B0(
        fu_LIFTING_n276), .Y(fu_LIFTING_n278) );
  AOI21X1 fu_LIFTING_U578 ( .A0(fu_LIFTING_n241), .A1(fu_LIFTING_n239), .B0(
        fu_LIFTING_n49), .Y(fu_LIFTING_n279) );
  AOI21X1 fu_LIFTING_U577 ( .A0(fu_LIFTING_n37), .A1(fu_LIFTING_N78), .B0(
        fu_LIFTING_n279), .Y(fu_LIFTING_n281) );
  AOI21X1 fu_LIFTING_U576 ( .A0(fu_LIFTING_n241), .A1(fu_LIFTING_n239), .B0(
        fu_LIFTING_n50), .Y(fu_LIFTING_n282) );
  AOI21X1 fu_LIFTING_U575 ( .A0(fu_LIFTING_n37), .A1(fu_LIFTING_N79), .B0(
        fu_LIFTING_n282), .Y(fu_LIFTING_n284) );
  AOI21X1 fu_LIFTING_U574 ( .A0(fu_LIFTING_n241), .A1(fu_LIFTING_n239), .B0(
        fu_LIFTING_n52), .Y(fu_LIFTING_n285) );
  AOI21X1 fu_LIFTING_U573 ( .A0(fu_LIFTING_n37), .A1(fu_LIFTING_N80), .B0(
        fu_LIFTING_n285), .Y(fu_LIFTING_n287) );
  AOI21X1 fu_LIFTING_U572 ( .A0(fu_LIFTING_n241), .A1(fu_LIFTING_n239), .B0(
        fu_LIFTING_n53), .Y(fu_LIFTING_n288) );
  AOI21X1 fu_LIFTING_U571 ( .A0(fu_LIFTING_n37), .A1(fu_LIFTING_N81), .B0(
        fu_LIFTING_n288), .Y(fu_LIFTING_n290) );
  AOI21X1 fu_LIFTING_U570 ( .A0(fu_LIFTING_n241), .A1(fu_LIFTING_n239), .B0(
        fu_LIFTING_n54), .Y(fu_LIFTING_n291) );
  AOI21X1 fu_LIFTING_U569 ( .A0(fu_LIFTING_n37), .A1(fu_LIFTING_N82), .B0(
        fu_LIFTING_n291), .Y(fu_LIFTING_n293) );
  AOI21X1 fu_LIFTING_U568 ( .A0(fu_LIFTING_n241), .A1(fu_LIFTING_n239), .B0(
        fu_LIFTING_n55), .Y(fu_LIFTING_n294) );
  AOI21X1 fu_LIFTING_U567 ( .A0(fu_LIFTING_n37), .A1(fu_LIFTING_N83), .B0(
        fu_LIFTING_n294), .Y(fu_LIFTING_n296) );
  AOI21X1 fu_LIFTING_U566 ( .A0(fu_LIFTING_n241), .A1(fu_LIFTING_n239), .B0(
        fu_LIFTING_n56), .Y(fu_LIFTING_n297) );
  AOI21X1 fu_LIFTING_U565 ( .A0(fu_LIFTING_n37), .A1(fu_LIFTING_N84), .B0(
        fu_LIFTING_n297), .Y(fu_LIFTING_n299) );
  AOI21X1 fu_LIFTING_U564 ( .A0(fu_LIFTING_n241), .A1(fu_LIFTING_n239), .B0(
        fu_LIFTING_n57), .Y(fu_LIFTING_n300) );
  AOI21X1 fu_LIFTING_U563 ( .A0(fu_LIFTING_n37), .A1(fu_LIFTING_N85), .B0(
        fu_LIFTING_n300), .Y(fu_LIFTING_n302) );
  AOI222X2 fu_LIFTING_U562 ( .A0(fu_LIFTING_N65), .A1(fu_LIFTING_n36), .B0(
        fu_LIFTING_n83), .B1(fu_LIFTING_N425), .C0(fu_LIFTING_n235), .C1(
        fu_LIFTING_N305), .Y(fu_LIFTING_n374) );
  AOI21X1 fu_LIFTING_U561 ( .A0(fu_LIFTING_n241), .A1(fu_LIFTING_n239), .B0(
        fu_LIFTING_n59), .Y(fu_LIFTING_n303) );
  AOI21X1 fu_LIFTING_U560 ( .A0(fu_LIFTING_n37), .A1(fu_LIFTING_N86), .B0(
        fu_LIFTING_n303), .Y(fu_LIFTING_n305) );
  AOI222X2 fu_LIFTING_U559 ( .A0(fu_LIFTING_N64), .A1(fu_LIFTING_n36), .B0(
        fu_LIFTING_n83), .B1(fu_LIFTING_N424), .C0(fu_LIFTING_n37), .C1(
        fu_LIFTING_N544), .Y(fu_LIFTING_n376) );
  AOI21X1 fu_LIFTING_U558 ( .A0(fu_LIFTING_n241), .A1(fu_LIFTING_n239), .B0(
        fu_LIFTING_n60), .Y(fu_LIFTING_n306) );
  AOI21X1 fu_LIFTING_U557 ( .A0(fu_LIFTING_n37), .A1(fu_LIFTING_N87), .B0(
        fu_LIFTING_n306), .Y(fu_LIFTING_n308) );
  AOI222X2 fu_LIFTING_U556 ( .A0(fu_LIFTING_N63), .A1(fu_LIFTING_n36), .B0(
        fu_LIFTING_n83), .B1(fu_LIFTING_N423), .C0(fu_LIFTING_n235), .C1(
        fu_LIFTING_N303), .Y(fu_LIFTING_n378) );
  AOI21X1 fu_LIFTING_U555 ( .A0(fu_LIFTING_n36), .A1(fu_LIFTING_N88), .B0(
        fu_LIFTING_n309), .Y(fu_LIFTING_n311) );
  AOI222X2 fu_LIFTING_U554 ( .A0(fu_LIFTING_N62), .A1(fu_LIFTING_n36), .B0(
        fu_LIFTING_n83), .B1(fu_LIFTING_N422), .C0(fu_LIFTING_n235), .C1(
        fu_LIFTING_N302), .Y(fu_LIFTING_n380) );
  AOI21X1 fu_LIFTING_U553 ( .A0(fu_LIFTING_n241), .A1(fu_LIFTING_n239), .B0(
        fu_LIFTING_n61), .Y(fu_LIFTING_n312) );
  AOI21X1 fu_LIFTING_U552 ( .A0(fu_LIFTING_n37), .A1(fu_LIFTING_N89), .B0(
        fu_LIFTING_n312), .Y(fu_LIFTING_n314) );
  AOI222X2 fu_LIFTING_U551 ( .A0(fu_LIFTING_N61), .A1(fu_LIFTING_n36), .B0(
        fu_LIFTING_n83), .B1(fu_LIFTING_N421), .C0(fu_LIFTING_n235), .C1(
        fu_LIFTING_N301), .Y(fu_LIFTING_n382) );
  AOI21X1 fu_LIFTING_U550 ( .A0(fu_LIFTING_n241), .A1(fu_LIFTING_n239), .B0(
        fu_LIFTING_n64), .Y(fu_LIFTING_n315) );
  AOI21X1 fu_LIFTING_U549 ( .A0(fu_LIFTING_n37), .A1(fu_LIFTING_N90), .B0(
        fu_LIFTING_n315), .Y(fu_LIFTING_n317) );
  AOI222X2 fu_LIFTING_U548 ( .A0(fu_LIFTING_N60), .A1(fu_LIFTING_n36), .B0(
        fu_LIFTING_n83), .B1(fu_LIFTING_N420), .C0(fu_LIFTING_n235), .C1(
        fu_LIFTING_N300), .Y(fu_LIFTING_n384) );
  AOI21X1 fu_LIFTING_U547 ( .A0(fu_LIFTING_n241), .A1(fu_LIFTING_n239), .B0(
        fu_LIFTING_n66), .Y(fu_LIFTING_n318) );
  AOI21X1 fu_LIFTING_U546 ( .A0(fu_LIFTING_n37), .A1(fu_LIFTING_N91), .B0(
        fu_LIFTING_n318), .Y(fu_LIFTING_n320) );
  AOI222X2 fu_LIFTING_U545 ( .A0(fu_LIFTING_N59), .A1(fu_LIFTING_n36), .B0(
        fu_LIFTING_n83), .B1(fu_LIFTING_N419), .C0(fu_LIFTING_n235), .C1(
        fu_LIFTING_N299), .Y(fu_LIFTING_n386) );
  AOI21X1 fu_LIFTING_U544 ( .A0(fu_LIFTING_n241), .A1(fu_LIFTING_n239), .B0(
        fu_LIFTING_n67), .Y(fu_LIFTING_n321) );
  AOI21X1 fu_LIFTING_U543 ( .A0(fu_LIFTING_n37), .A1(fu_LIFTING_N92), .B0(
        fu_LIFTING_n321), .Y(fu_LIFTING_n323) );
  AOI222X2 fu_LIFTING_U542 ( .A0(fu_LIFTING_N58), .A1(fu_LIFTING_n36), .B0(
        fu_LIFTING_n83), .B1(fu_LIFTING_N418), .C0(fu_LIFTING_n235), .C1(
        fu_LIFTING_N298), .Y(fu_LIFTING_n388) );
  AOI21X1 fu_LIFTING_U541 ( .A0(fu_LIFTING_n408), .A1(fu_LIFTING_N93), .B0(
        fu_LIFTING_n324), .Y(fu_LIFTING_n326) );
  AOI222X2 fu_LIFTING_U540 ( .A0(fu_LIFTING_N57), .A1(fu_LIFTING_n36), .B0(
        fu_LIFTING_n83), .B1(fu_LIFTING_N417), .C0(fu_LIFTING_n235), .C1(
        fu_LIFTING_N297), .Y(fu_LIFTING_n390) );
  AOI21X1 fu_LIFTING_U539 ( .A0(fu_LIFTING_n241), .A1(fu_LIFTING_n239), .B0(
        fu_LIFTING_n71), .Y(fu_LIFTING_n327) );
  AOI21X1 fu_LIFTING_U538 ( .A0(fu_LIFTING_n37), .A1(fu_LIFTING_N94), .B0(
        fu_LIFTING_n327), .Y(fu_LIFTING_n329) );
  AOI222X2 fu_LIFTING_U537 ( .A0(fu_LIFTING_N56), .A1(fu_LIFTING_n36), .B0(
        fu_LIFTING_n83), .B1(fu_LIFTING_N416), .C0(fu_LIFTING_n235), .C1(
        fu_LIFTING_N296), .Y(fu_LIFTING_n392) );
  AOI21X1 fu_LIFTING_U536 ( .A0(fu_LIFTING_n241), .A1(fu_LIFTING_n239), .B0(
        fu_LIFTING_n81), .Y(fu_LIFTING_n330) );
  AOI21X1 fu_LIFTING_U535 ( .A0(fu_LIFTING_n37), .A1(fu_LIFTING_N95), .B0(
        fu_LIFTING_n330), .Y(fu_LIFTING_n332) );
  AOI222X2 fu_LIFTING_U534 ( .A0(fu_LIFTING_N55), .A1(fu_LIFTING_n36), .B0(
        fu_LIFTING_n83), .B1(fu_LIFTING_N415), .C0(fu_LIFTING_n235), .C1(
        fu_LIFTING_N295), .Y(fu_LIFTING_n394) );
  AOI21X1 fu_LIFTING_U533 ( .A0(fu_LIFTING_n241), .A1(fu_LIFTING_n239), .B0(
        fu_LIFTING_n82), .Y(fu_LIFTING_n333) );
  AOI21X1 fu_LIFTING_U532 ( .A0(fu_LIFTING_n37), .A1(fu_LIFTING_N96), .B0(
        fu_LIFTING_n333), .Y(fu_LIFTING_n335) );
  AOI222X2 fu_LIFTING_U531 ( .A0(fu_LIFTING_N54), .A1(fu_LIFTING_n36), .B0(
        fu_LIFTING_n83), .B1(fu_LIFTING_N414), .C0(fu_LIFTING_n235), .C1(
        fu_LIFTING_N294), .Y(fu_LIFTING_n396) );
  AOI21X1 fu_LIFTING_U530 ( .A0(fu_LIFTING_n236), .A1(fu_LIFTING_n237), .B0(
        fu_LIFTING_n79), .Y(fu_LIFTING_n336) );
  AOI21X1 fu_LIFTING_U529 ( .A0(fu_LIFTING_n83), .A1(fu_LIFTING_N697), .B0(
        fu_LIFTING_n336), .Y(fu_LIFTING_n338) );
  AOI222X2 fu_LIFTING_U528 ( .A0(fu_LIFTING_N53), .A1(fu_LIFTING_n36), .B0(
        fu_LIFTING_n83), .B1(fu_LIFTING_N413), .C0(fu_LIFTING_n235), .C1(
        fu_LIFTING_N293), .Y(fu_LIFTING_n398) );
  AOI21X1 fu_LIFTING_U527 ( .A0(fu_LIFTING_n36), .A1(fu_LIFTING_N98), .B0(
        fu_LIFTING_n340), .Y(fu_LIFTING_n342) );
  AOI21X1 fu_LIFTING_U526 ( .A0(fu_LIFTING_n241), .A1(fu_LIFTING_n239), .B0(
        fu_LIFTING_n343), .Y(fu_LIFTING_n344) );
  AOI21X1 fu_LIFTING_U525 ( .A0(fu_LIFTING_n37), .A1(fu_LIFTING_N99), .B0(
        fu_LIFTING_n344), .Y(fu_LIFTING_n346) );
  AOI21X1 fu_LIFTING_U524 ( .A0(fu_LIFTING_n241), .A1(fu_LIFTING_n239), .B0(
        fu_LIFTING_n350), .Y(fu_LIFTING_n347) );
  AOI21X1 fu_LIFTING_U523 ( .A0(fu_LIFTING_n37), .A1(fu_LIFTING_N644), .B0(
        fu_LIFTING_n347), .Y(fu_LIFTING_n349) );
  AOI21X1 fu_LIFTING_U522 ( .A0(fu_LIFTING_n36), .A1(fu_LIFTING_N645), .B0(
        fu_LIFTING_n351), .Y(fu_LIFTING_n353) );
  AOI21X1 fu_LIFTING_U521 ( .A0(fu_LIFTING_n236), .A1(fu_LIFTING_n237), .B0(
        fu_LIFTING_n40), .Y(fu_LIFTING_n355) );
  AOI21X1 fu_LIFTING_U520 ( .A0(fu_LIFTING_n83), .A1(fu_LIFTING_N702), .B0(
        fu_LIFTING_n355), .Y(fu_LIFTING_n357) );
  AOI21X1 fu_LIFTING_U519 ( .A0(fu_LIFTING_n241), .A1(fu_LIFTING_n239), .B0(
        fu_LIFTING_n70), .Y(fu_LIFTING_n358) );
  AOI21X1 fu_LIFTING_U518 ( .A0(fu_LIFTING_n37), .A1(fu_LIFTING_N647), .B0(
        fu_LIFTING_n358), .Y(fu_LIFTING_n360) );
  AOI21X1 fu_LIFTING_U517 ( .A0(fu_LIFTING_n241), .A1(fu_LIFTING_n239), .B0(
        fu_LIFTING_n262), .Y(fu_LIFTING_n254) );
  AOI21X1 fu_LIFTING_U516 ( .A0(fu_LIFTING_n37), .A1(fu_LIFTING_N72), .B0(
        fu_LIFTING_n254), .Y(fu_LIFTING_n261) );
  CLKMX2X12 fu_LIFTING_U515 ( .A(fu_LIFTING_reg_x1_23_), .B(
        rf_RF_t1data_wire[23]), .S0(fu_LIFTING_n249), .Y(fu_LIFTING_N80) );
  CLKMX2X12 fu_LIFTING_U514 ( .A(fu_LIFTING_reg_x1_22_), .B(
        rf_RF_t1data_wire[22]), .S0(fu_LIFTING_n249), .Y(fu_LIFTING_N81) );
  CLKMX2X12 fu_LIFTING_U513 ( .A(fu_LIFTING_reg_x1_21_), .B(
        rf_RF_t1data_wire[21]), .S0(fu_LIFTING_n249), .Y(fu_LIFTING_N82) );
  CLKMX2X12 fu_LIFTING_U512 ( .A(fu_LIFTING_reg_x1_20_), .B(
        rf_RF_t1data_wire[20]), .S0(fu_LIFTING_n249), .Y(fu_LIFTING_N83) );
  CLKMX2X12 fu_LIFTING_U511 ( .A(fu_LIFTING_reg_x1_19_), .B(
        rf_RF_t1data_wire[19]), .S0(fu_LIFTING_n249), .Y(fu_LIFTING_N84) );
  CLKMX2X12 fu_LIFTING_U510 ( .A(fu_LIFTING_reg_x1_17_), .B(
        rf_RF_t1data_wire[17]), .S0(fu_LIFTING_n42), .Y(fu_LIFTING_N86) );
  CLKMX2X12 fu_LIFTING_U509 ( .A(fu_LIFTING_reg_x1_16_), .B(
        rf_RF_t1data_wire[16]), .S0(fu_LIFTING_n42), .Y(fu_LIFTING_N87) );
  CLKMX2X12 fu_LIFTING_U508 ( .A(fu_LIFTING_reg_x1_12_), .B(n1820), .S0(
        fu_LIFTING_n42), .Y(fu_LIFTING_N91) );
  OAI211X2 fu_LIFTING_U507 ( .A0(fu_LIFTING_n266), .A1(fu_LIFTING_n1), .B0(
        fu_LIFTING_n265), .C0(fu_LIFTING_n264), .Y(fu_LIFTING_n473) );
  OAI21X1 fu_LIFTING_U506 ( .A0(fu_LIFTING_n36), .A1(fu_LIFTING_n234), .B0(
        fu_LIFTING_N78), .Y(fu_LIFTING_n280) );
  OAI21X1 fu_LIFTING_U505 ( .A0(fu_LIFTING_n36), .A1(fu_LIFTING_n234), .B0(
        fu_LIFTING_N80), .Y(fu_LIFTING_n286) );
  OAI21X1 fu_LIFTING_U504 ( .A0(fu_LIFTING_n36), .A1(fu_LIFTING_n234), .B0(
        fu_LIFTING_N81), .Y(fu_LIFTING_n289) );
  OAI21X1 fu_LIFTING_U503 ( .A0(fu_LIFTING_n36), .A1(fu_LIFTING_n234), .B0(
        fu_LIFTING_N82), .Y(fu_LIFTING_n292) );
  OAI21X1 fu_LIFTING_U502 ( .A0(fu_LIFTING_n36), .A1(fu_LIFTING_n234), .B0(
        fu_LIFTING_N83), .Y(fu_LIFTING_n295) );
  AOI222X2 fu_LIFTING_U501 ( .A0(fu_LIFTING_N667), .A1(fu_LIFTING_n240), .B0(
        fu_LIFTING_n37), .B1(fu_LIFTING_N547), .C0(fu_LIFTING_n238), .C1(
        fu_LIFTING_N187), .Y(fu_LIFTING_n369) );
  OAI21X1 fu_LIFTING_U500 ( .A0(fu_LIFTING_n36), .A1(fu_LIFTING_n234), .B0(
        fu_LIFTING_N84), .Y(fu_LIFTING_n298) );
  AOI222X2 fu_LIFTING_U499 ( .A0(fu_LIFTING_N666), .A1(fu_LIFTING_n240), .B0(
        fu_LIFTING_n37), .B1(fu_LIFTING_N546), .C0(fu_LIFTING_n238), .C1(
        fu_LIFTING_N186), .Y(fu_LIFTING_n371) );
  AOI222X2 fu_LIFTING_U498 ( .A0(fu_LIFTING_N665), .A1(fu_LIFTING_n240), .B0(
        fu_LIFTING_n37), .B1(fu_LIFTING_N545), .C0(fu_LIFTING_n238), .C1(
        fu_LIFTING_N185), .Y(fu_LIFTING_n373) );
  OAI21X1 fu_LIFTING_U497 ( .A0(fu_LIFTING_n36), .A1(fu_LIFTING_n234), .B0(
        fu_LIFTING_N86), .Y(fu_LIFTING_n304) );
  AOI222X2 fu_LIFTING_U496 ( .A0(fu_LIFTING_N664), .A1(fu_LIFTING_n240), .B0(
        fu_LIFTING_n234), .B1(fu_LIFTING_N304), .C0(fu_LIFTING_n238), .C1(
        fu_LIFTING_N184), .Y(fu_LIFTING_n375) );
  OAI21X1 fu_LIFTING_U495 ( .A0(fu_LIFTING_n36), .A1(fu_LIFTING_n233), .B0(
        fu_LIFTING_N87), .Y(fu_LIFTING_n307) );
  AOI222X2 fu_LIFTING_U494 ( .A0(fu_LIFTING_N663), .A1(fu_LIFTING_n240), .B0(
        fu_LIFTING_n37), .B1(fu_LIFTING_N543), .C0(fu_LIFTING_n475), .C1(
        fu_LIFTING_N183), .Y(fu_LIFTING_n377) );
  AOI222X2 fu_LIFTING_U493 ( .A0(fu_LIFTING_N662), .A1(fu_LIFTING_n240), .B0(
        fu_LIFTING_n37), .B1(fu_LIFTING_N542), .C0(fu_LIFTING_n475), .C1(
        fu_LIFTING_N182), .Y(fu_LIFTING_n379) );
  OAI21X1 fu_LIFTING_U492 ( .A0(fu_LIFTING_n36), .A1(fu_LIFTING_n233), .B0(
        fu_LIFTING_N89), .Y(fu_LIFTING_n313) );
  AOI222X2 fu_LIFTING_U491 ( .A0(fu_LIFTING_N661), .A1(fu_LIFTING_n240), .B0(
        fu_LIFTING_n37), .B1(fu_LIFTING_N541), .C0(fu_LIFTING_n475), .C1(
        fu_LIFTING_N181), .Y(fu_LIFTING_n381) );
  AOI222X2 fu_LIFTING_U490 ( .A0(fu_LIFTING_N660), .A1(fu_LIFTING_n240), .B0(
        fu_LIFTING_n37), .B1(fu_LIFTING_N540), .C0(fu_LIFTING_n238), .C1(
        fu_LIFTING_N180), .Y(fu_LIFTING_n383) );
  OAI21X1 fu_LIFTING_U489 ( .A0(fu_LIFTING_n36), .A1(fu_LIFTING_n233), .B0(
        fu_LIFTING_N91), .Y(fu_LIFTING_n319) );
  AOI222X2 fu_LIFTING_U488 ( .A0(fu_LIFTING_N659), .A1(fu_LIFTING_n476), .B0(
        fu_LIFTING_n37), .B1(fu_LIFTING_N539), .C0(fu_LIFTING_n238), .C1(
        fu_LIFTING_N179), .Y(fu_LIFTING_n385) );
  OAI21X1 fu_LIFTING_U487 ( .A0(fu_LIFTING_n36), .A1(fu_LIFTING_n233), .B0(
        fu_LIFTING_N92), .Y(fu_LIFTING_n322) );
  AOI222X2 fu_LIFTING_U486 ( .A0(fu_LIFTING_N658), .A1(fu_LIFTING_n476), .B0(
        fu_LIFTING_n37), .B1(fu_LIFTING_N538), .C0(fu_LIFTING_n238), .C1(
        fu_LIFTING_N178), .Y(fu_LIFTING_n387) );
  AOI222X2 fu_LIFTING_U485 ( .A0(fu_LIFTING_N657), .A1(fu_LIFTING_n240), .B0(
        fu_LIFTING_n37), .B1(fu_LIFTING_N537), .C0(fu_LIFTING_n238), .C1(
        fu_LIFTING_N177), .Y(fu_LIFTING_n389) );
  OAI21X1 fu_LIFTING_U484 ( .A0(fu_LIFTING_n36), .A1(fu_LIFTING_n233), .B0(
        fu_LIFTING_N94), .Y(fu_LIFTING_n328) );
  AOI222X2 fu_LIFTING_U483 ( .A0(fu_LIFTING_N656), .A1(fu_LIFTING_n240), .B0(
        fu_LIFTING_n37), .B1(fu_LIFTING_N536), .C0(fu_LIFTING_n238), .C1(
        fu_LIFTING_N176), .Y(fu_LIFTING_n391) );
  OAI21X1 fu_LIFTING_U482 ( .A0(fu_LIFTING_n36), .A1(fu_LIFTING_n233), .B0(
        fu_LIFTING_N95), .Y(fu_LIFTING_n331) );
  OAI21X1 fu_LIFTING_U481 ( .A0(fu_LIFTING_n36), .A1(fu_LIFTING_n233), .B0(
        fu_LIFTING_N96), .Y(fu_LIFTING_n334) );
  OAI21X1 fu_LIFTING_U480 ( .A0(fu_LIFTING_n36), .A1(fu_LIFTING_n233), .B0(
        fu_LIFTING_N644), .Y(fu_LIFTING_n348) );
  OAI21X1 fu_LIFTING_U479 ( .A0(fu_LIFTING_n36), .A1(fu_LIFTING_n234), .B0(
        fu_LIFTING_N647), .Y(fu_LIFTING_n359) );
  AOI222X2 fu_LIFTING_U478 ( .A0(fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_28_), 
        .A1(fu_LIFTING_n242), .B0(fu_LIFTING_n243), .B1(
        fu_LIFTING_reg_out_tmp_28_), .C0(fu_LIFTING_n246), .C1(
        ic_socket_LIFTING_o1_data0_wire[28]), .Y(fu_LIFTING_n439) );
  AOI222X2 fu_LIFTING_U477 ( .A0(fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_27_), 
        .A1(fu_LIFTING_n242), .B0(fu_LIFTING_n243), .B1(
        fu_LIFTING_reg_out_tmp_27_), .C0(fu_LIFTING_n246), .C1(
        ic_socket_LIFTING_o1_data0_wire[27]), .Y(fu_LIFTING_n438) );
  AOI222X2 fu_LIFTING_U476 ( .A0(fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_26_), 
        .A1(fu_LIFTING_n242), .B0(fu_LIFTING_n243), .B1(
        fu_LIFTING_reg_out_tmp_26_), .C0(fu_LIFTING_n247), .C1(
        ic_socket_LIFTING_o1_data0_wire[26]), .Y(fu_LIFTING_n437) );
  AOI222X2 fu_LIFTING_U475 ( .A0(fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_25_), 
        .A1(fu_LIFTING_n242), .B0(fu_LIFTING_n243), .B1(
        fu_LIFTING_reg_out_tmp_25_), .C0(fu_LIFTING_n247), .C1(
        ic_socket_LIFTING_o1_data0_wire[25]), .Y(fu_LIFTING_n436) );
  AOI222X2 fu_LIFTING_U474 ( .A0(fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_24_), 
        .A1(fu_LIFTING_n242), .B0(fu_LIFTING_n243), .B1(
        fu_LIFTING_reg_out_tmp_24_), .C0(fu_LIFTING_n247), .C1(
        ic_socket_LIFTING_o1_data0_wire[24]), .Y(fu_LIFTING_n435) );
  AOI222X2 fu_LIFTING_U473 ( .A0(fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_23_), 
        .A1(fu_LIFTING_n242), .B0(fu_LIFTING_n243), .B1(
        fu_LIFTING_reg_out_tmp_23_), .C0(fu_LIFTING_n247), .C1(
        ic_socket_LIFTING_o1_data0_wire[23]), .Y(fu_LIFTING_n434) );
  AOI222X2 fu_LIFTING_U472 ( .A0(fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_22_), 
        .A1(fu_LIFTING_n242), .B0(fu_LIFTING_n243), .B1(
        fu_LIFTING_reg_out_tmp_22_), .C0(fu_LIFTING_n247), .C1(
        ic_socket_LIFTING_o1_data0_wire[22]), .Y(fu_LIFTING_n433) );
  AOI222X2 fu_LIFTING_U471 ( .A0(fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_21_), 
        .A1(fu_LIFTING_n242), .B0(fu_LIFTING_n243), .B1(
        fu_LIFTING_reg_out_tmp_21_), .C0(fu_LIFTING_n247), .C1(
        ic_socket_LIFTING_o1_data0_wire[21]), .Y(fu_LIFTING_n432) );
  AOI222X2 fu_LIFTING_U470 ( .A0(fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_20_), 
        .A1(fu_LIFTING_n242), .B0(fu_LIFTING_n243), .B1(
        fu_LIFTING_reg_out_tmp_20_), .C0(fu_LIFTING_n246), .C1(
        ic_socket_LIFTING_o1_data0_wire[20]), .Y(fu_LIFTING_n431) );
  AOI222X2 fu_LIFTING_U469 ( .A0(fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_19_), 
        .A1(fu_LIFTING_n242), .B0(fu_LIFTING_n243), .B1(
        fu_LIFTING_reg_out_tmp_19_), .C0(fu_LIFTING_n246), .C1(
        ic_socket_LIFTING_o1_data0_wire[19]), .Y(fu_LIFTING_n430) );
  AOI222X2 fu_LIFTING_U468 ( .A0(fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_18_), 
        .A1(fu_LIFTING_n242), .B0(fu_LIFTING_n243), .B1(
        fu_LIFTING_reg_out_tmp_18_), .C0(fu_LIFTING_n246), .C1(
        ic_socket_LIFTING_o1_data0_wire[18]), .Y(fu_LIFTING_n429) );
  AOI222X2 fu_LIFTING_U467 ( .A0(fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_17_), 
        .A1(fu_LIFTING_n242), .B0(fu_LIFTING_n243), .B1(
        fu_LIFTING_reg_out_tmp_17_), .C0(fu_LIFTING_n246), .C1(
        ic_socket_LIFTING_o1_data0_wire[17]), .Y(fu_LIFTING_n428) );
  AOI222X2 fu_LIFTING_U466 ( .A0(fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_16_), 
        .A1(fu_LIFTING_n242), .B0(fu_LIFTING_n243), .B1(
        fu_LIFTING_reg_out_tmp_16_), .C0(fu_LIFTING_n246), .C1(
        ic_socket_LIFTING_o1_data0_wire[16]), .Y(fu_LIFTING_n427) );
  AOI222X2 fu_LIFTING_U465 ( .A0(fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_15_), 
        .A1(fu_LIFTING_n242), .B0(fu_LIFTING_n243), .B1(
        fu_LIFTING_reg_out_tmp_15_), .C0(fu_LIFTING_n246), .C1(
        ic_socket_LIFTING_o1_data0_wire[15]), .Y(fu_LIFTING_n426) );
  AOI222X2 fu_LIFTING_U464 ( .A0(fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_14_), 
        .A1(fu_LIFTING_n242), .B0(fu_LIFTING_n243), .B1(
        fu_LIFTING_reg_out_tmp_14_), .C0(fu_LIFTING_n246), .C1(
        ic_socket_LIFTING_o1_data0_wire[14]), .Y(fu_LIFTING_n425) );
  AOI222X2 fu_LIFTING_U463 ( .A0(fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_13_), 
        .A1(fu_LIFTING_n242), .B0(fu_LIFTING_n243), .B1(
        fu_LIFTING_reg_out_tmp_13_), .C0(fu_LIFTING_n246), .C1(
        ic_socket_LIFTING_o1_data0_wire[13]), .Y(fu_LIFTING_n424) );
  AOI222X2 fu_LIFTING_U462 ( .A0(fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_12_), 
        .A1(fu_LIFTING_n242), .B0(fu_LIFTING_n243), .B1(
        fu_LIFTING_reg_out_tmp_12_), .C0(fu_LIFTING_n246), .C1(
        ic_socket_LIFTING_o1_data0_wire[12]), .Y(fu_LIFTING_n423) );
  OR2X2 fu_LIFTING_U461 ( .A(fu_LIFTING_t1opcode_wire[1]), .B(
        fu_LIFTING_t1opcode_wire[2]), .Y(fu_LIFTING_n251) );
  NAND2BX2 fu_LIFTING_U460 ( .AN(fu_LIFTING_n72), .B(
        fu_LIFTING_t1opcode_wire[2]), .Y(fu_LIFTING_n255) );
  NAND2BX2 fu_LIFTING_U459 ( .AN(fu_LIFTING_n72), .B(
        fu_LIFTING_t1opcode_wire[1]), .Y(fu_LIFTING_n259) );
  AOI21X1 fu_LIFTING_U458 ( .A0(fu_LIFTING_n37), .A1(fu_LIFTING_N74), .B0(
        fu_LIFTING_n267), .Y(fu_LIFTING_n269) );
  OAI211X2 fu_LIFTING_U457 ( .A0(fu_LIFTING_n43), .A1(fu_LIFTING_n1), .B0(
        fu_LIFTING_n269), .C0(fu_LIFTING_n268), .Y(fu_LIFTING_n472) );
  OAI211X2 fu_LIFTING_U456 ( .A0(fu_LIFTING_n44), .A1(fu_LIFTING_n1), .B0(
        fu_LIFTING_n272), .C0(fu_LIFTING_n271), .Y(fu_LIFTING_n471) );
  AOI22X1 fu_LIFTING_U455 ( .A0(fu_LIFTING_n238), .A1(fu_LIFTING_N677), .B0(
        fu_LIFTING_N77), .B1(fu_LIFTING_n234), .Y(fu_LIFTING_n277) );
  AOI22X1 fu_LIFTING_U454 ( .A0(fu_LIFTING_n83), .A1(fu_LIFTING_N679), .B0(
        fu_LIFTING_N79), .B1(fu_LIFTING_n234), .Y(fu_LIFTING_n283) );
  CLKMX2X12 fu_LIFTING_U453 ( .A(fu_LIFTING_reg_x1_11_), .B(
        rf_RF_t1data_wire[11]), .S0(fu_LIFTING_n42), .Y(fu_LIFTING_N92) );
  NAND2X2 fu_LIFTING_U452 ( .A(fu_LIFTING_n384), .B(fu_LIFTING_n383), .Y(
        fu_LIFTING_n489) );
  AOI222X4 fu_LIFTING_U451 ( .A0(fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_31_), 
        .A1(fu_LIFTING_n242), .B0(fu_LIFTING_n243), .B1(
        fu_LIFTING_reg_out_tmp_31_), .C0(fu_LIFTING_n246), .C1(
        ic_socket_LIFTING_o1_data0_wire[31]), .Y(fu_LIFTING_n442) );
  CLKMX2X12 fu_LIFTING_U450 ( .A(fu_LIFTING_reg_x1_9_), .B(n1812), .S0(
        fu_LIFTING_n42), .Y(fu_LIFTING_N94) );
  AOI222X2 fu_LIFTING_U449 ( .A0(fu_LIFTING_N66), .A1(fu_LIFTING_n36), .B0(
        fu_LIFTING_n83), .B1(fu_LIFTING_N426), .C0(fu_LIFTING_n235), .C1(
        fu_LIFTING_N306), .Y(fu_LIFTING_n372) );
  NAND2X2 fu_LIFTING_U448 ( .A(fu_LIFTING_n402), .B(fu_LIFTING_n401), .Y(
        fu_LIFTING_n480) );
  AOI222X4 fu_LIFTING_U447 ( .A0(fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_30_), 
        .A1(fu_LIFTING_n242), .B0(fu_LIFTING_n243), .B1(
        fu_LIFTING_reg_out_tmp_30_), .C0(fu_LIFTING_n246), .C1(
        ic_socket_LIFTING_o1_data0_wire[30]), .Y(fu_LIFTING_n441) );
  NAND2X8 fu_LIFTING_U446 ( .A(fu_LIFTING_n362), .B(fu_LIFTING_n361), .Y(
        fu_LIFTING_n500) );
  MX2X8 fu_LIFTING_U445 ( .A(fu_LIFTING_reg_x2_0_), .B(n2111), .S0(
        fu_LIFTING_n248), .Y(fu_LIFTING_N703) );
  ADDFX1 fu_LIFTING_U444 ( .A(fu_LIFTING_mult_96_DP_OP_281_6650_6_n74), .B(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n75), .CI(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n23), .CO(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n22), .S(fu_LIFTING_N650) );
  ADDFX1 fu_LIFTING_U443 ( .A(fu_LIFTING_mult_96_DP_OP_281_6650_6_n72), .B(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n73), .CI(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n22), .CO(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n21), .S(fu_LIFTING_N651) );
  ADDFX1 fu_LIFTING_U442 ( .A(fu_LIFTING_mult_96_DP_OP_281_6650_6_n54), .B(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n55), .CI(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n13), .CO(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n12), .S(fu_LIFTING_N660) );
  ADDFX1 fu_LIFTING_U441 ( .A(fu_LIFTING_mult_96_DP_OP_281_6650_6_n52), .B(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n53), .CI(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n12), .CO(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n11), .S(fu_LIFTING_N661) );
  ADDFX1 fu_LIFTING_U440 ( .A(fu_LIFTING_mult_96_DP_OP_281_6650_6_n50), .B(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n51), .CI(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n11), .CO(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n10), .S(fu_LIFTING_N662) );
  OAI2BB1X4 fu_LIFTING_U439 ( .A0N(fu_LIFTING_N647), .A1N(fu_LIFTING_n135), 
        .B0(fu_LIFTING_n134), .Y(fu_LIFTING_mult_96_DP_OP_281_6650_6_n25) );
  AOI222X4 fu_LIFTING_U438 ( .A0(fu_LIFTING_N98), .A1(fu_LIFTING_n133), .B0(
        fu_LIFTING_N98), .B1(fu_LIFTING_n39), .C0(fu_LIFTING_n133), .C1(
        fu_LIFTING_n39), .Y(fu_LIFTING_n135) );
  AOI222X4 fu_LIFTING_U437 ( .A0(fu_LIFTING_N646), .A1(fu_LIFTING_n78), .B0(
        fu_LIFTING_N646), .B1(fu_LIFTING_n132), .C0(fu_LIFTING_n78), .C1(
        fu_LIFTING_n132), .Y(fu_LIFTING_n133) );
  XOR3X4 fu_LIFTING_U436 ( .A(fu_LIFTING_n131), .B(fu_LIFTING_n130), .C(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n33), .Y(fu_LIFTING_N671) );
  ADDFX1 fu_LIFTING_U435 ( .A(fu_LIFTING_mult_92_DP_OP_280_6650_5_n66), .B(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n67), .CI(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n19), .CO(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n18), .S(fu_LIFTING_N534) );
  ADDFX1 fu_LIFTING_U434 ( .A(fu_LIFTING_mult_92_DP_OP_280_6650_5_n56), .B(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n57), .CI(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n14), .CO(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n13), .S(fu_LIFTING_N539) );
  ADDFX1 fu_LIFTING_U433 ( .A(fu_LIFTING_mult_92_DP_OP_280_6650_5_n50), .B(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n51), .CI(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n11), .CO(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n10), .S(fu_LIFTING_N542) );
  ADDFX1 fu_LIFTING_U432 ( .A(fu_LIFTING_mult_92_DP_OP_280_6650_5_n48), .B(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n49), .CI(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n10), .CO(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n9), .S(fu_LIFTING_N543) );
  ADDFX1 fu_LIFTING_U431 ( .A(fu_LIFTING_mult_92_DP_OP_280_6650_5_n46), .B(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n47), .CI(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n9), .CO(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n8), .S(fu_LIFTING_N544) );
  ADDFX1 fu_LIFTING_U430 ( .A(fu_LIFTING_mult_92_DP_OP_280_6650_5_n44), .B(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n45), .CI(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n8), .CO(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n7), .S(fu_LIFTING_N545) );
  ADDFX2 fu_LIFTING_U429 ( .A(fu_LIFTING_mult_92_DP_OP_280_6650_5_n36), .B(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n37), .CI(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n4), .CO(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n3), .S(fu_LIFTING_N549) );
  CLKXOR2X4 fu_LIFTING_U428 ( .A(fu_LIFTING_N673), .B(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n2), .Y(fu_LIFTING_n122) );
  OAI2BB1X4 fu_LIFTING_U427 ( .A0N(fu_LIFTING_N703), .A1N(fu_LIFTING_n127), 
        .B0(fu_LIFTING_n126), .Y(fu_LIFTING_n129) );
  AOI222X4 fu_LIFTING_U426 ( .A0(fu_LIFTING_N699), .A1(fu_LIFTING_n125), .B0(
        fu_LIFTING_N699), .B1(fu_LIFTING_n76), .C0(fu_LIFTING_n125), .C1(
        fu_LIFTING_n76), .Y(fu_LIFTING_n127) );
  OAI21BX4 fu_LIFTING_U425 ( .A0(fu_LIFTING_N703), .A1(fu_LIFTING_n124), .B0N(
        fu_LIFTING_N700), .Y(fu_LIFTING_n125) );
  XNOR2X2 fu_LIFTING_U424 ( .A(fu_LIFTING_N73), .B(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n2), .Y(fu_LIFTING_n117) );
  OA21X4 fu_LIFTING_U423 ( .A0(fu_LIFTING_mult_88_DP_OP_277_6650_4_n81), .A1(
        fu_LIFTING_N644), .B0(fu_LIFTING_N647), .Y(fu_LIFTING_n119) );
  ADDFX1 fu_LIFTING_U422 ( .A(fu_LIFTING_mult_88_DP_OP_277_6650_4_n53), .B(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n54), .CI(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n14), .CO(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n13), .S(fu_LIFTING_N419) );
  ADDFX1 fu_LIFTING_U421 ( .A(fu_LIFTING_mult_88_DP_OP_277_6650_4_n43), .B(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n44), .CI(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n9), .CO(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n8), .S(fu_LIFTING_N424) );
  OAI2BB1X2 fu_LIFTING_U420 ( .A0N(fu_LIFTING_mult_88_DP_OP_277_6650_4_n78), 
        .A1N(fu_LIFTING_n121), .B0(fu_LIFTING_n120), .Y(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n25) );
  ADDFX1 fu_LIFTING_U419 ( .A(fu_LIFTING_mult_84_DP_OP_276_6650_3_n74), .B(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n75), .CI(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n24), .CO(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n23), .S(fu_LIFTING_N289) );
  ADDFX1 fu_LIFTING_U418 ( .A(fu_LIFTING_mult_84_DP_OP_276_6650_3_n72), .B(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n73), .CI(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n23), .CO(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n22), .S(fu_LIFTING_N290) );
  ADDFX1 fu_LIFTING_U417 ( .A(fu_LIFTING_mult_84_DP_OP_276_6650_3_n60), .B(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n61), .CI(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n17), .CO(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n16), .S(fu_LIFTING_N296) );
  ADDFX1 fu_LIFTING_U416 ( .A(fu_LIFTING_mult_84_DP_OP_276_6650_3_n58), .B(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n59), .CI(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n16), .CO(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n15), .S(fu_LIFTING_N297) );
  ADDFX1 fu_LIFTING_U415 ( .A(fu_LIFTING_mult_84_DP_OP_276_6650_3_n56), .B(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n57), .CI(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n15), .CO(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n14), .S(fu_LIFTING_N298) );
  ADDFX1 fu_LIFTING_U414 ( .A(fu_LIFTING_mult_84_DP_OP_276_6650_3_n54), .B(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n55), .CI(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n14), .CO(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n13), .S(fu_LIFTING_N299) );
  ADDFX1 fu_LIFTING_U413 ( .A(fu_LIFTING_mult_84_DP_OP_276_6650_3_n42), .B(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n43), .CI(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n8), .CO(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n7), .S(fu_LIFTING_N305) );
  ADDFX2 fu_LIFTING_U412 ( .A(fu_LIFTING_mult_84_DP_OP_276_6650_3_n36), .B(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n37), .CI(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n5), .CO(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n4), .S(fu_LIFTING_N308) );
  ADDFX2 fu_LIFTING_U411 ( .A(fu_LIFTING_mult_84_DP_OP_276_6650_3_n34), .B(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n35), .CI(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n4), .CO(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n3), .S(fu_LIFTING_N309) );
  OAI21X4 fu_LIFTING_U410 ( .A0(fu_LIFTING_mult_84_DP_OP_276_6650_3_n79), .A1(
        fu_LIFTING_n115), .B0(fu_LIFTING_mult_84_DP_OP_276_6650_3_n78), .Y(
        fu_LIFTING_n114) );
  OAI21X2 fu_LIFTING_U409 ( .A0(fu_LIFTING_mult_84_DP_OP_276_6650_3_n83), .A1(
        fu_LIFTING_n111), .B0(fu_LIFTING_mult_84_DP_OP_276_6650_3_n82), .Y(
        fu_LIFTING_n110) );
  OA21X4 fu_LIFTING_U408 ( .A0(fu_LIFTING_mult_84_DP_OP_276_6650_3_n84), .A1(
        fu_LIFTING_N700), .B0(fu_LIFTING_N703), .Y(fu_LIFTING_n111) );
  OAI2BB1X4 fu_LIFTING_U407 ( .A0N(fu_LIFTING_mult_84_DP_OP_276_6650_3_n79), 
        .A1N(fu_LIFTING_n115), .B0(fu_LIFTING_n114), .Y(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n25) );
  OAI2BB1X4 fu_LIFTING_U406 ( .A0N(fu_LIFTING_mult_84_DP_OP_276_6650_3_n81), 
        .A1N(fu_LIFTING_n113), .B0(fu_LIFTING_n112), .Y(fu_LIFTING_n115) );
  OAI2BB1X4 fu_LIFTING_U405 ( .A0N(fu_LIFTING_mult_84_DP_OP_276_6650_3_n83), 
        .A1N(fu_LIFTING_n111), .B0(fu_LIFTING_n110), .Y(fu_LIFTING_n113) );
  XNOR2X4 fu_LIFTING_U404 ( .A(fu_LIFTING_N672), .B(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n2), .Y(fu_LIFTING_n109) );
  ADDFX2 fu_LIFTING_U403 ( .A(fu_LIFTING_mult_79_DP_OP_279_6650_2_n62), .B(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n63), .CI(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n19), .CO(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n18), .S(fu_LIFTING_N174) );
  OA21X4 fu_LIFTING_U402 ( .A0(fu_LIFTING_mult_79_DP_OP_279_6650_2_n78), .A1(
        fu_LIFTING_N99), .B0(fu_LIFTING_N647), .Y(fu_LIFTING_n106) );
  ADDFX1 fu_LIFTING_U401 ( .A(fu_LIFTING_mult_79_DP_OP_279_6650_2_n52), .B(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n53), .CI(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n14), .CO(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n13), .S(fu_LIFTING_N179) );
  ADDFX1 fu_LIFTING_U400 ( .A(fu_LIFTING_mult_79_DP_OP_279_6650_2_n44), .B(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n45), .CI(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n10), .CO(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n9), .S(fu_LIFTING_N183) );
  ADDFX1 fu_LIFTING_U399 ( .A(fu_LIFTING_mult_79_DP_OP_279_6650_2_n42), .B(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n43), .CI(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n9), .CO(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n8), .S(fu_LIFTING_N184) );
  OAI2BB1X1 fu_LIFTING_U398 ( .A0N(fu_LIFTING_mult_79_DP_OP_279_6650_2_n77), 
        .A1N(fu_LIFTING_n106), .B0(fu_LIFTING_n105), .Y(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n25) );
  OAI21X1 fu_LIFTING_U397 ( .A0(fu_LIFTING_mult_79_DP_OP_279_6650_2_n77), .A1(
        fu_LIFTING_n106), .B0(fu_LIFTING_mult_79_DP_OP_279_6650_2_n76), .Y(
        fu_LIFTING_n105) );
  ADDFHX4 fu_LIFTING_U396 ( .A(fu_LIFTING_mult_75_DP_OP_278_6650_1_n65), .B(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n67), .CI(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n12), .CO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n11), .S(fu_LIFTING_N61) );
  ADDFX2 fu_LIFTING_U395 ( .A(fu_LIFTING_mult_75_DP_OP_278_6650_1_n92), .B(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n94), .CI(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n21), .CO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n20), .S(fu_LIFTING_N52) );
  ADDFX1 fu_LIFTING_U394 ( .A(fu_LIFTING_mult_75_DP_OP_278_6650_1_n89), .B(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n91), .CI(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n20), .CO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n19), .S(fu_LIFTING_N53) );
  ADDFX1 fu_LIFTING_U393 ( .A(fu_LIFTING_mult_75_DP_OP_278_6650_1_n74), .B(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n76), .CI(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n15), .CO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n14), .S(fu_LIFTING_N58) );
  ADDFX1 fu_LIFTING_U392 ( .A(fu_LIFTING_mult_75_DP_OP_278_6650_1_n71), .B(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n73), .CI(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n14), .CO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n13), .S(fu_LIFTING_N59) );
  ADDFX1 fu_LIFTING_U391 ( .A(fu_LIFTING_mult_75_DP_OP_278_6650_1_n62), .B(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n64), .CI(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n11), .CO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n10), .S(fu_LIFTING_N62) );
  AND3X2 fu_LIFTING_U390 ( .A(fu_LIFTING_N700), .B(fu_LIFTING_N702), .C(
        fu_LIFTING_N703), .Y(fu_LIFTING_n94) );
  INVX4 fu_LIFTING_U389 ( .A(fu_LIFTING_mult_75_DP_OP_278_6650_1_n116), .Y(
        fu_LIFTING_n95) );
  OAI2BB1X4 fu_LIFTING_U388 ( .A0N(fu_LIFTING_mult_75_DP_OP_278_6650_1_n114), 
        .A1N(fu_LIFTING_n98), .B0(fu_LIFTING_n97), .Y(fu_LIFTING_n100) );
  AOI222X4 fu_LIFTING_U387 ( .A0(fu_LIFTING_n96), .A1(fu_LIFTING_n70), .B0(
        fu_LIFTING_n96), .B1(fu_LIFTING_n95), .C0(fu_LIFTING_n70), .C1(
        fu_LIFTING_n95), .Y(fu_LIFTING_n98) );
  OAI2BB1X4 fu_LIFTING_U386 ( .A0N(fu_LIFTING_mult_75_DP_OP_278_6650_1_n111), 
        .A1N(fu_LIFTING_n100), .B0(fu_LIFTING_n99), .Y(fu_LIFTING_n102) );
  OAI22X4 fu_LIFTING_U385 ( .A0(fu_LIFTING_n94), .A1(fu_LIFTING_N701), .B0(
        fu_LIFTING_N700), .B1(fu_LIFTING_N702), .Y(fu_LIFTING_n96) );
  XOR2X8 fu_LIFTING_U384 ( .A(fu_LIFTING_n41), .B(fu_LIFTING_n500), .Y(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n47) );
  ADDFHX4 fu_LIFTING_U383 ( .A(fu_LIFTING_sub_98_DP_OP_282_1544_7_n47), .B(
        fu_LIFTING_n466), .CI(fu_LIFTING_sub_98_DP_OP_282_1544_7_n10), .CO(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n9), .S(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_23_) );
  ADDFHX4 fu_LIFTING_U382 ( .A(fu_LIFTING_sub_98_DP_OP_282_1544_7_n40), .B(
        fu_LIFTING_n473), .CI(fu_LIFTING_sub_98_DP_OP_282_1544_7_n3), .CO(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n2), .S(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_30_) );
  XOR2X8 fu_LIFTING_U381 ( .A(fu_LIFTING_sub_98_DP_OP_282_1544_7_n2), .B(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n1), .Y(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_31_) );
  CLKXOR2X2 fu_LIFTING_U380 ( .A(fu_LIFTING_n41), .B(fu_LIFTING_n492), .Y(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n55) );
  CLKXOR2X2 fu_LIFTING_U379 ( .A(fu_LIFTING_n41), .B(fu_LIFTING_n491), .Y(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n56) );
  CLKBUFX24 fu_LIFTING_U378 ( .A(fu_LIFTING_n74), .Y(fu_LIFTING_n243) );
  CLKMX2X12 fu_LIFTING_U377 ( .A(fu_LIFTING_reg_x1_5_), .B(
        rf_RF_t1data_wire[5]), .S0(fu_LIFTING_n42), .Y(fu_LIFTING_N98) );
  ADDHX2 fu_LIFTING_U376 ( .A(fu_LIFTING_N98), .B(fu_LIFTING_N646), .CO(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n77), .S(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n78) );
  CLKMX2X12 fu_LIFTING_U375 ( .A(fu_LIFTING_reg_x2_4_), .B(n1825), .S0(
        fu_LIFTING_n248), .Y(fu_LIFTING_N699) );
  ADDFX2 fu_LIFTING_U374 ( .A(fu_LIFTING_N699), .B(fu_LIFTING_N698), .CI(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n115), .CO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n111), .S(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n112) );
  ADDHX2 fu_LIFTING_U373 ( .A(fu_LIFTING_N699), .B(fu_LIFTING_N700), .CO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n115), .S(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n116) );
  ADDHX2 fu_LIFTING_U372 ( .A(fu_LIFTING_N699), .B(fu_LIFTING_N702), .CO(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n83), .S(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n84) );
  NAND2BX8 fu_LIFTING_U371 ( .AN(fu_LIFTING_n247), .B(rstx), .Y(fu_LIFTING_n72) );
  NOR2BX8 fu_LIFTING_U370 ( .AN(fu_LIFTING_n107), .B(fu_LIFTING_n72), .Y(
        fu_LIFTING_N993) );
  AOI222X2 fu_LIFTING_U369 ( .A0(fu_LIFTING_N652), .A1(fu_LIFTING_n240), .B0(
        fu_LIFTING_n37), .B1(fu_LIFTING_N532), .C0(fu_LIFTING_n238), .C1(
        fu_LIFTING_N172), .Y(fu_LIFTING_n399) );
  AOI222X2 fu_LIFTING_U368 ( .A0(fu_LIFTING_N649), .A1(fu_LIFTING_n240), .B0(
        fu_LIFTING_n234), .B1(fu_LIFTING_N289), .C0(fu_LIFTING_n238), .C1(
        fu_LIFTING_N169), .Y(fu_LIFTING_n405) );
  CLKINVX32 fu_LIFTING_U367 ( .A(fu_LIFTING_n240), .Y(fu_LIFTING_n241) );
  NOR2X2 fu_LIFTING_U366 ( .A(fu_LIFTING_N702), .B(fu_LIFTING_N701), .Y(
        fu_LIFTING_n124) );
  NAND2X2 fu_LIFTING_U365 ( .A(fu_LIFTING_n88), .B(fu_LIFTING_n89), .Y(
        fu_LIFTING_n132) );
  ADDFX4 fu_LIFTING_U364 ( .A(fu_LIFTING_sub_98_DP_OP_282_1544_7_n46), .B(
        fu_LIFTING_n467), .CI(fu_LIFTING_sub_98_DP_OP_282_1544_7_n9), .CO(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n8), .S(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_24_) );
  ADDHX2 fu_LIFTING_U363 ( .A(fu_LIFTING_N99), .B(fu_LIFTING_N646), .CO(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n80), .S(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n81) );
  OAI21X1 fu_LIFTING_U362 ( .A0(fu_LIFTING_mult_88_DP_OP_277_6650_4_n80), .A1(
        fu_LIFTING_n119), .B0(fu_LIFTING_mult_88_DP_OP_277_6650_4_n79), .Y(
        fu_LIFTING_n118) );
  OAI2BB1X2 fu_LIFTING_U361 ( .A0N(fu_LIFTING_mult_88_DP_OP_277_6650_4_n80), 
        .A1N(fu_LIFTING_n119), .B0(fu_LIFTING_n118), .Y(fu_LIFTING_n121) );
  XNOR2X2 fu_LIFTING_U360 ( .A(fu_LIFTING_N676), .B(fu_LIFTING_N677), .Y(
        fu_LIFTING_n90) );
  XNOR2X2 fu_LIFTING_U359 ( .A(fu_LIFTING_N78), .B(fu_LIFTING_N77), .Y(
        fu_LIFTING_n103) );
  XOR3X2 fu_LIFTING_U358 ( .A(fu_LIFTING_mult_79_DP_OP_279_6650_2_n29), .B(
        fu_LIFTING_n104), .C(fu_LIFTING_n103), .Y(fu_LIFTING_N191) );
  ADDFX1 fu_LIFTING_U357 ( .A(fu_LIFTING_mult_92_DP_OP_280_6650_5_n74), .B(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n75), .CI(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n23), .CO(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n22), .S(fu_LIFTING_N530) );
  ADDFX1 fu_LIFTING_U356 ( .A(fu_LIFTING_mult_84_DP_OP_276_6650_3_n70), .B(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n71), .CI(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n22), .CO(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n21), .S(fu_LIFTING_N291) );
  ADDFX1 fu_LIFTING_U355 ( .A(fu_LIFTING_mult_88_DP_OP_277_6650_4_n67), .B(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n68), .CI(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n21), .CO(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n20), .S(fu_LIFTING_N412) );
  ADDFX1 fu_LIFTING_U354 ( .A(fu_LIFTING_mult_79_DP_OP_279_6650_2_n60), .B(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n61), .CI(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n18), .CO(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n17), .S(fu_LIFTING_N175) );
  ADDFX1 fu_LIFTING_U353 ( .A(fu_LIFTING_mult_84_DP_OP_276_6650_3_n52), .B(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n53), .CI(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n13), .CO(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n12), .S(fu_LIFTING_N300) );
  ADDFX1 fu_LIFTING_U352 ( .A(fu_LIFTING_mult_88_DP_OP_277_6650_4_n49), .B(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n50), .CI(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n12), .CO(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n11), .S(fu_LIFTING_N421) );
  CLKBUFX24 fu_LIFTING_U351 ( .A(n2211), .Y(fu_LIFTING_n246) );
  INVX20 fu_LIFTING_U350 ( .A(fu_LIFTING_n238), .Y(fu_LIFTING_n239) );
  CLKMX2X12 fu_LIFTING_U349 ( .A(fu_LIFTING_reg_x1_8_), .B(
        rf_RF_t1data_wire[8]), .S0(fu_LIFTING_n42), .Y(fu_LIFTING_N95) );
  CLKMX2X12 fu_LIFTING_U348 ( .A(fu_LIFTING_reg_x1_7_), .B(n1814), .S0(
        fu_LIFTING_n42), .Y(fu_LIFTING_N96) );
  ADDFX1 fu_LIFTING_U347 ( .A(fu_LIFTING_N96), .B(fu_LIFTING_N92), .CI(
        fu_LIFTING_N95), .CO(fu_LIFTING_mult_88_DP_OP_277_6650_4_n66), .S(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n67) );
  ADDFX1 fu_LIFTING_U346 ( .A(fu_LIFTING_N97), .B(fu_LIFTING_N93), .CI(
        fu_LIFTING_N96), .CO(fu_LIFTING_mult_88_DP_OP_277_6650_4_n68), .S(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n69) );
  INVX12 fu_LIFTING_U345 ( .A(n1757), .Y(fu_LIFTING_n249) );
  CLKXOR2X2 fu_LIFTING_U344 ( .A(fu_LIFTING_n41), .B(fu_LIFTING_n484), .Y(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n63) );
  OAI2BB1X2 fu_LIFTING_U343 ( .A0N(fu_LIFTING_n87), .A1N(fu_LIFTING_n102), 
        .B0(fu_LIFTING_n101), .Y(fu_LIFTING_mult_75_DP_OP_278_6650_1_n25) );
  BUFX2 fu_LIFTING_U342 ( .A(fu_LIFTING_mult_75_DP_OP_278_6650_1_n109), .Y(
        fu_LIFTING_n87) );
  ADDHX2 fu_LIFTING_U341 ( .A(fu_LIFTING_n73), .B(fu_LIFTING_N701), .CO(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n81), .S(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n82) );
  OAI2BB1X2 fu_LIFTING_U340 ( .A0N(fu_LIFTING_mult_92_DP_OP_280_6650_5_n81), 
        .A1N(fu_LIFTING_n129), .B0(fu_LIFTING_n128), .Y(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n25) );
  OAI21X1 fu_LIFTING_U339 ( .A0(fu_LIFTING_mult_92_DP_OP_280_6650_5_n81), .A1(
        fu_LIFTING_n129), .B0(fu_LIFTING_mult_92_DP_OP_280_6650_5_n80), .Y(
        fu_LIFTING_n128) );
  CMPR42X2 fu_LIFTING_U338 ( .A(fu_LIFTING_N687), .B(fu_LIFTING_N688), .C(
        fu_LIFTING_N684), .D(fu_LIFTING_N683), .ICI(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n69), .S(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n68), .ICO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n66), .CO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n67) );
  OAI211X2 fu_LIFTING_U337 ( .A0(fu_LIFTING_n49), .A1(fu_LIFTING_n1), .B0(
        fu_LIFTING_n281), .C0(fu_LIFTING_n280), .Y(fu_LIFTING_n468) );
  OAI211X2 fu_LIFTING_U336 ( .A0(fu_LIFTING_n52), .A1(fu_LIFTING_n1), .B0(
        fu_LIFTING_n287), .C0(fu_LIFTING_n286), .Y(fu_LIFTING_n466) );
  ADDFX2 fu_LIFTING_U335 ( .A(fu_LIFTING_mult_92_DP_OP_280_6650_5_n72), .B(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n73), .CI(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n22), .CO(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n21), .S(fu_LIFTING_N531) );
  CLKBUFX24 fu_LIFTING_U334 ( .A(fu_LIFTING_n75), .Y(fu_LIFTING_n242) );
  AOI222X2 fu_LIFTING_U333 ( .A0(fu_LIFTING_N291), .A1(fu_LIFTING_n234), .B0(
        fu_LIFTING_n83), .B1(fu_LIFTING_N411), .C0(fu_LIFTING_n238), .C1(
        fu_LIFTING_N171), .Y(fu_LIFTING_n401) );
  NOR3X8 fu_LIFTING_U332 ( .A(fu_LIFTING_n72), .B(fu_LIFTING_n252), .C(
        fu_LIFTING_n251), .Y(fu_LIFTING_n476) );
  NOR2X4 fu_LIFTING_U331 ( .A(fu_LIFTING_n259), .B(fu_LIFTING_n258), .Y(
        fu_LIFTING_n407) );
  BUFX12 fu_LIFTING_U330 ( .A(fu_LIFTING_n407), .Y(fu_LIFTING_n233) );
  ADDHX4 fu_LIFTING_U329 ( .A(fu_LIFTING_N702), .B(fu_LIFTING_N703), .CO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n113), .S(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n114) );
  OAI21X4 fu_LIFTING_U328 ( .A0(fu_LIFTING_mult_75_DP_OP_278_6650_1_n114), 
        .A1(fu_LIFTING_n98), .B0(fu_LIFTING_mult_75_DP_OP_278_6650_1_n112), 
        .Y(fu_LIFTING_n97) );
  CLKXOR2X2 fu_LIFTING_U327 ( .A(fu_LIFTING_n41), .B(fu_LIFTING_n481), .Y(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n66) );
  XNOR2X2 fu_LIFTING_U326 ( .A(fu_LIFTING_N77), .B(fu_LIFTING_N76), .Y(
        fu_LIFTING_n116) );
  XNOR2X2 fu_LIFTING_U325 ( .A(fu_LIFTING_N676), .B(fu_LIFTING_N675), .Y(
        fu_LIFTING_n108) );
  OAI21X1 fu_LIFTING_U324 ( .A0(fu_LIFTING_N647), .A1(fu_LIFTING_n135), .B0(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n80), .Y(fu_LIFTING_n134) );
  NAND2BX2 fu_LIFTING_U323 ( .AN(fu_LIFTING_t1opcode_wire[2]), .B(
        fu_LIFTING_t1opcode_wire[0]), .Y(fu_LIFTING_n250) );
  INVX2 fu_LIFTING_U322 ( .A(fu_LIFTING_t1opcode_wire[0]), .Y(fu_LIFTING_n252)
         );
  OR2X2 fu_LIFTING_U321 ( .A(fu_LIFTING_t1opcode_wire[2]), .B(
        fu_LIFTING_t1opcode_wire[0]), .Y(fu_LIFTING_n258) );
  NOR2X2 fu_LIFTING_U320 ( .A(fu_LIFTING_t1opcode_wire[1]), .B(
        fu_LIFTING_t1opcode_wire[0]), .Y(fu_LIFTING_n256) );
  NAND2BX2 fu_LIFTING_U319 ( .AN(fu_LIFTING_t1opcode_wire[1]), .B(
        fu_LIFTING_t1opcode_wire[0]), .Y(fu_LIFTING_n253) );
  NOR2X6 fu_LIFTING_U318 ( .A(fu_LIFTING_n246), .B(fu_LIFTING_n107), .Y(
        fu_LIFTING_n74) );
  AOI21X6 fu_LIFTING_U317 ( .A0(fu_LIFTING_t1opcode_wire[2]), .A1(
        fu_LIFTING_t1opcode_wire[1]), .B0(fu_LIFTING_n246), .Y(fu_LIFTING_n75)
         );
  NOR2BX4 fu_LIFTING_U316 ( .AN(fu_LIFTING_n248), .B(fu_LIFTING_n72), .Y(
        fu_LIFTING_N929) );
  CLKBUFX24 fu_LIFTING_U315 ( .A(fu_LIFTING_N961), .Y(fu_LIFTING_n85) );
  OR3X2 fu_LIFTING_U314 ( .A(fu_LIFTING_n72), .B(fu_LIFTING_t1opcode_wire[0]), 
        .C(fu_LIFTING_n251), .Y(fu_LIFTING_n231) );
  CLKBUFX24 fu_LIFTING_U313 ( .A(fu_LIFTING_N993), .Y(fu_LIFTING_n84) );
  INVX2 fu_LIFTING_U312 ( .A(fu_LIFTING_n255), .Y(fu_LIFTING_n257) );
  NOR2X6 fu_LIFTING_U311 ( .A(fu_LIFTING_n255), .B(fu_LIFTING_n253), .Y(
        fu_LIFTING_n475) );
  BUFX20 fu_LIFTING_U310 ( .A(fu_LIFTING_n476), .Y(fu_LIFTING_n240) );
  BUFX14 fu_LIFTING_U309 ( .A(fu_LIFTING_N929), .Y(fu_LIFTING_n245) );
  BUFX14 fu_LIFTING_U308 ( .A(fu_LIFTING_N929), .Y(fu_LIFTING_n244) );
  CLKBUFX20 fu_LIFTING_U307 ( .A(fu_LIFTING_n407), .Y(fu_LIFTING_n234) );
  CLKBUFX32 fu_LIFTING_U306 ( .A(fu_LIFTING_n475), .Y(fu_LIFTING_n238) );
  AND2X2 fu_LIFTING_U305 ( .A(fu_LIFTING_n257), .B(fu_LIFTING_n256), .Y(
        fu_LIFTING_n408) );
  BUFX14 fu_LIFTING_U304 ( .A(fu_LIFTING_n233), .Y(fu_LIFTING_n235) );
  INVX4 fu_LIFTING_U303 ( .A(fu_LIFTING_N696), .Y(fu_LIFTING_n82) );
  INVX4 fu_LIFTING_U302 ( .A(fu_LIFTING_N695), .Y(fu_LIFTING_n81) );
  INVX2 fu_LIFTING_U301 ( .A(fu_LIFTING_N697), .Y(fu_LIFTING_n80) );
  INVX2 fu_LIFTING_U300 ( .A(fu_LIFTING_N97), .Y(fu_LIFTING_n79) );
  INVX4 fu_LIFTING_U299 ( .A(fu_LIFTING_N99), .Y(fu_LIFTING_n78) );
  INVX2 fu_LIFTING_U298 ( .A(fu_LIFTING_N644), .Y(fu_LIFTING_n77) );
  INVX2 fu_LIFTING_U297 ( .A(fu_LIFTING_N96), .Y(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n104) );
  INVX2 fu_LIFTING_U296 ( .A(fu_LIFTING_N95), .Y(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n103) );
  INVX2 fu_LIFTING_U295 ( .A(fu_LIFTING_N700), .Y(fu_LIFTING_n350) );
  INVX4 fu_LIFTING_U294 ( .A(fu_LIFTING_N702), .Y(fu_LIFTING_n76) );
  AOI22X2 fu_LIFTING_U293 ( .A0(fu_LIFTING_n238), .A1(fu_LIFTING_N697), .B0(
        fu_LIFTING_N97), .B1(fu_LIFTING_n233), .Y(fu_LIFTING_n337) );
  AOI22X2 fu_LIFTING_U292 ( .A0(fu_LIFTING_n83), .A1(fu_LIFTING_N699), .B0(
        fu_LIFTING_N99), .B1(fu_LIFTING_n234), .Y(fu_LIFTING_n345) );
  INVX2 fu_LIFTING_U291 ( .A(fu_LIFTING_N699), .Y(fu_LIFTING_n343) );
  MX2X8 fu_LIFTING_U290 ( .A(fu_LIFTING_reg_x2_2_), .B(n1810), .S0(
        fu_LIFTING_n248), .Y(fu_LIFTING_N701) );
  INVX4 fu_LIFTING_U289 ( .A(fu_LIFTING_N698), .Y(fu_LIFTING_n73) );
  INVX2 fu_LIFTING_U288 ( .A(fu_LIFTING_N701), .Y(fu_LIFTING_n354) );
  AOI22X2 fu_LIFTING_U287 ( .A0(fu_LIFTING_n238), .A1(fu_LIFTING_N701), .B0(
        fu_LIFTING_N645), .B1(fu_LIFTING_n233), .Y(fu_LIFTING_n352) );
  AOI22X2 fu_LIFTING_U286 ( .A0(fu_LIFTING_n238), .A1(fu_LIFTING_N702), .B0(
        fu_LIFTING_N646), .B1(fu_LIFTING_n233), .Y(fu_LIFTING_n356) );
  INVX4 fu_LIFTING_U285 ( .A(fu_LIFTING_N694), .Y(fu_LIFTING_n71) );
  AOI22X2 fu_LIFTING_U284 ( .A0(fu_LIFTING_n238), .A1(fu_LIFTING_N698), .B0(
        fu_LIFTING_N98), .B1(fu_LIFTING_n233), .Y(fu_LIFTING_n341) );
  INVX2 fu_LIFTING_U283 ( .A(fu_LIFTING_N98), .Y(fu_LIFTING_n339) );
  ADDFX2 fu_LIFTING_U282 ( .A(fu_LIFTING_N646), .B(fu_LIFTING_N98), .CI(
        fu_LIFTING_N645), .CO(fu_LIFTING_mult_88_DP_OP_277_6650_4_n78), .S(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n79) );
  INVX2 fu_LIFTING_U281 ( .A(fu_LIFTING_N93), .Y(fu_LIFTING_n69) );
  INVX2 fu_LIFTING_U280 ( .A(fu_LIFTING_N94), .Y(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n102) );
  INVX4 fu_LIFTING_U279 ( .A(fu_LIFTING_N693), .Y(fu_LIFTING_n68) );
  AOI22X2 fu_LIFTING_U278 ( .A0(fu_LIFTING_n238), .A1(fu_LIFTING_N693), .B0(
        fu_LIFTING_N93), .B1(fu_LIFTING_n234), .Y(fu_LIFTING_n325) );
  OAI211X2 fu_LIFTING_U277 ( .A0(fu_LIFTING_n350), .A1(fu_LIFTING_n2), .B0(
        fu_LIFTING_n349), .C0(fu_LIFTING_n348), .Y(fu_LIFTING_n446) );
  INVX4 fu_LIFTING_U276 ( .A(fu_LIFTING_N692), .Y(fu_LIFTING_n67) );
  OAI211X2 fu_LIFTING_U275 ( .A0(fu_LIFTING_n354), .A1(fu_LIFTING_n241), .B0(
        fu_LIFTING_n353), .C0(fu_LIFTING_n352), .Y(fu_LIFTING_n445) );
  INVX4 fu_LIFTING_U274 ( .A(fu_LIFTING_N691), .Y(fu_LIFTING_n66) );
  INVX2 fu_LIFTING_U273 ( .A(fu_LIFTING_N91), .Y(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n99) );
  INVX2 fu_LIFTING_U272 ( .A(fu_LIFTING_N92), .Y(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n100) );
  INVX4 fu_LIFTING_U271 ( .A(fu_LIFTING_N688), .Y(fu_LIFTING_n63) );
  AOI22X2 fu_LIFTING_U270 ( .A0(fu_LIFTING_n83), .A1(fu_LIFTING_N690), .B0(
        fu_LIFTING_N90), .B1(fu_LIFTING_n234), .Y(fu_LIFTING_n316) );
  INVX4 fu_LIFTING_U269 ( .A(fu_LIFTING_N689), .Y(fu_LIFTING_n61) );
  AOI22X2 fu_LIFTING_U268 ( .A0(fu_LIFTING_n238), .A1(fu_LIFTING_N688), .B0(
        fu_LIFTING_N88), .B1(fu_LIFTING_n234), .Y(fu_LIFTING_n310) );
  INVX4 fu_LIFTING_U267 ( .A(fu_LIFTING_N687), .Y(fu_LIFTING_n60) );
  INVX2 fu_LIFTING_U266 ( .A(fu_LIFTING_N89), .Y(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n97) );
  INVX2 fu_LIFTING_U265 ( .A(fu_LIFTING_N87), .Y(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n95) );
  INVX4 fu_LIFTING_U264 ( .A(fu_LIFTING_N686), .Y(fu_LIFTING_n59) );
  INVX2 fu_LIFTING_U263 ( .A(fu_LIFTING_N86), .Y(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n94) );
  INVX4 fu_LIFTING_U262 ( .A(fu_LIFTING_N684), .Y(fu_LIFTING_n56) );
  AOI22X2 fu_LIFTING_U261 ( .A0(fu_LIFTING_n83), .A1(fu_LIFTING_N685), .B0(
        fu_LIFTING_N85), .B1(fu_LIFTING_n234), .Y(fu_LIFTING_n301) );
  INVX4 fu_LIFTING_U260 ( .A(fu_LIFTING_N683), .Y(fu_LIFTING_n55) );
  INVX2 fu_LIFTING_U259 ( .A(fu_LIFTING_N84), .Y(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n92) );
  INVX2 fu_LIFTING_U258 ( .A(fu_LIFTING_N83), .Y(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n91) );
  INVX4 fu_LIFTING_U257 ( .A(fu_LIFTING_N682), .Y(fu_LIFTING_n54) );
  AOI222X2 fu_LIFTING_U256 ( .A0(fu_LIFTING_N648), .A1(fu_LIFTING_n240), .B0(
        fu_LIFTING_n83), .B1(fu_LIFTING_N408), .C0(fu_LIFTING_n37), .C1(
        fu_LIFTING_N528), .Y(fu_LIFTING_n409) );
  INVX4 fu_LIFTING_U255 ( .A(fu_LIFTING_N681), .Y(fu_LIFTING_n53) );
  INVX2 fu_LIFTING_U254 ( .A(fu_LIFTING_N82), .Y(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n90) );
  NAND2X2 fu_LIFTING_U253 ( .A(fu_LIFTING_n410), .B(fu_LIFTING_n409), .Y(
        fu_LIFTING_n477) );
  AOI222X2 fu_LIFTING_U252 ( .A0(fu_LIFTING_N49), .A1(fu_LIFTING_n36), .B0(
        fu_LIFTING_n83), .B1(fu_LIFTING_N409), .C0(fu_LIFTING_n37), .C1(
        fu_LIFTING_N529), .Y(fu_LIFTING_n406) );
  INVX2 fu_LIFTING_U251 ( .A(fu_LIFTING_N81), .Y(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n89) );
  INVX4 fu_LIFTING_U250 ( .A(fu_LIFTING_N79), .Y(fu_LIFTING_n51) );
  CLKXOR2X2 fu_LIFTING_U249 ( .A(fu_LIFTING_n41), .B(fu_LIFTING_n477), .Y(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n70) );
  NAND2X2 fu_LIFTING_U248 ( .A(fu_LIFTING_n406), .B(fu_LIFTING_n405), .Y(
        fu_LIFTING_n478) );
  AOI222X2 fu_LIFTING_U247 ( .A0(fu_LIFTING_N50), .A1(fu_LIFTING_n36), .B0(
        fu_LIFTING_n83), .B1(fu_LIFTING_N410), .C0(fu_LIFTING_n37), .C1(
        fu_LIFTING_N530), .Y(fu_LIFTING_n404) );
  AOI222X2 fu_LIFTING_U246 ( .A0(fu_LIFTING_N51), .A1(fu_LIFTING_n36), .B0(
        fu_LIFTING_n37), .B1(fu_LIFTING_N531), .C0(fu_LIFTING_n240), .C1(
        fu_LIFTING_N651), .Y(fu_LIFTING_n402) );
  CLKXOR2X2 fu_LIFTING_U245 ( .A(fu_LIFTING_n41), .B(fu_LIFTING_n478), .Y(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n69) );
  NAND2X2 fu_LIFTING_U244 ( .A(fu_LIFTING_n404), .B(fu_LIFTING_n403), .Y(
        fu_LIFTING_n479) );
  AOI222X2 fu_LIFTING_U243 ( .A0(fu_LIFTING_N653), .A1(fu_LIFTING_n240), .B0(
        fu_LIFTING_n37), .B1(fu_LIFTING_N533), .C0(fu_LIFTING_n238), .C1(
        fu_LIFTING_N173), .Y(fu_LIFTING_n397) );
  AOI222X2 fu_LIFTING_U242 ( .A0(fu_LIFTING_N52), .A1(fu_LIFTING_n36), .B0(
        fu_LIFTING_n83), .B1(fu_LIFTING_N412), .C0(fu_LIFTING_n235), .C1(
        fu_LIFTING_N292), .Y(fu_LIFTING_n400) );
  INVX2 fu_LIFTING_U241 ( .A(fu_LIFTING_N77), .Y(fu_LIFTING_n48) );
  AOI222X2 fu_LIFTING_U240 ( .A0(fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_0_), 
        .A1(fu_LIFTING_n242), .B0(fu_LIFTING_n243), .B1(
        fu_LIFTING_reg_out_tmp_0_), .C0(fu_LIFTING_n246), .C1(
        ic_socket_LIFTING_o1_data0_wire[0]), .Y(fu_LIFTING_n411) );
  INVX4 fu_LIFTING_U239 ( .A(fu_LIFTING_N677), .Y(fu_LIFTING_n47) );
  INVX2 fu_LIFTING_U238 ( .A(fu_LIFTING_N78), .Y(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n86) );
  AOI222X2 fu_LIFTING_U237 ( .A0(fu_LIFTING_N654), .A1(fu_LIFTING_n240), .B0(
        fu_LIFTING_n37), .B1(fu_LIFTING_N534), .C0(fu_LIFTING_n238), .C1(
        fu_LIFTING_N174), .Y(fu_LIFTING_n395) );
  INVX4 fu_LIFTING_U236 ( .A(fu_LIFTING_N76), .Y(fu_LIFTING_n45) );
  NAND2X2 fu_LIFTING_U235 ( .A(fu_LIFTING_n400), .B(fu_LIFTING_n399), .Y(
        fu_LIFTING_n481) );
  AOI222X2 fu_LIFTING_U234 ( .A0(fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_1_), 
        .A1(fu_LIFTING_n242), .B0(fu_LIFTING_n243), .B1(
        fu_LIFTING_reg_out_tmp_1_), .C0(fu_LIFTING_n246), .C1(
        ic_socket_LIFTING_o1_data0_wire[1]), .Y(fu_LIFTING_n412) );
  NAND2X2 fu_LIFTING_U233 ( .A(fu_LIFTING_n398), .B(fu_LIFTING_n397), .Y(
        fu_LIFTING_n482) );
  AOI22X2 fu_LIFTING_U232 ( .A0(fu_LIFTING_n238), .A1(fu_LIFTING_N676), .B0(
        fu_LIFTING_N76), .B1(fu_LIFTING_n233), .Y(fu_LIFTING_n274) );
  INVX4 fu_LIFTING_U231 ( .A(fu_LIFTING_N675), .Y(fu_LIFTING_n44) );
  AOI222X2 fu_LIFTING_U230 ( .A0(fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_2_), 
        .A1(fu_LIFTING_n75), .B0(fu_LIFTING_n243), .B1(
        fu_LIFTING_reg_out_tmp_2_), .C0(fu_LIFTING_n246), .C1(
        ic_socket_LIFTING_o1_data0_wire[2]), .Y(fu_LIFTING_n413) );
  AOI222X2 fu_LIFTING_U229 ( .A0(fu_LIFTING_N655), .A1(fu_LIFTING_n240), .B0(
        fu_LIFTING_n37), .B1(fu_LIFTING_N535), .C0(fu_LIFTING_n238), .C1(
        fu_LIFTING_N175), .Y(fu_LIFTING_n393) );
  AOI222X2 fu_LIFTING_U228 ( .A0(fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_3_), 
        .A1(fu_LIFTING_n242), .B0(fu_LIFTING_n243), .B1(
        fu_LIFTING_reg_out_tmp_3_), .C0(fu_LIFTING_n246), .C1(
        ic_socket_LIFTING_o1_data0_wire[3]), .Y(fu_LIFTING_n414) );
  INVX2 fu_LIFTING_U227 ( .A(fu_LIFTING_N75), .Y(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n83) );
  NAND2X2 fu_LIFTING_U226 ( .A(fu_LIFTING_n396), .B(fu_LIFTING_n395), .Y(
        fu_LIFTING_n483) );
  CLKXOR2X2 fu_LIFTING_U225 ( .A(fu_LIFTING_n41), .B(fu_LIFTING_n482), .Y(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n65) );
  NAND2X2 fu_LIFTING_U224 ( .A(fu_LIFTING_n394), .B(fu_LIFTING_n393), .Y(
        fu_LIFTING_n484) );
  CLKXOR2X2 fu_LIFTING_U223 ( .A(fu_LIFTING_n41), .B(fu_LIFTING_n483), .Y(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n64) );
  AOI222X2 fu_LIFTING_U222 ( .A0(fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_4_), 
        .A1(fu_LIFTING_n242), .B0(fu_LIFTING_n243), .B1(
        fu_LIFTING_reg_out_tmp_4_), .C0(fu_LIFTING_n246), .C1(
        ic_socket_LIFTING_o1_data0_wire[4]), .Y(fu_LIFTING_n415) );
  INVX4 fu_LIFTING_U221 ( .A(fu_LIFTING_N674), .Y(fu_LIFTING_n43) );
  AOI222X2 fu_LIFTING_U220 ( .A0(fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_5_), 
        .A1(fu_LIFTING_n242), .B0(fu_LIFTING_n74), .B1(
        fu_LIFTING_reg_out_tmp_5_), .C0(fu_LIFTING_n246), .C1(
        ic_socket_LIFTING_o1_data0_wire[5]), .Y(fu_LIFTING_n416) );
  MX2X4 fu_LIFTING_U219 ( .A(fu_LIFTING_reg_x2_30_), .B(n1862), .S0(
        fu_LIFTING_n248), .Y(fu_LIFTING_N673) );
  MX2X4 fu_LIFTING_U218 ( .A(fu_LIFTING_reg_x1_30_), .B(n1862), .S0(
        fu_LIFTING_n249), .Y(fu_LIFTING_N73) );
  MX2X4 fu_LIFTING_U217 ( .A(fu_LIFTING_reg_x2_31_), .B(n1860), .S0(
        fu_LIFTING_n248), .Y(fu_LIFTING_N672) );
  NAND2X2 fu_LIFTING_U216 ( .A(fu_LIFTING_n392), .B(fu_LIFTING_n391), .Y(
        fu_LIFTING_n485) );
  MX2X2 fu_LIFTING_U215 ( .A(fu_LIFTING_reg_x1_31_), .B(n1860), .S0(
        fu_LIFTING_n249), .Y(fu_LIFTING_N72) );
  INVX2 fu_LIFTING_U214 ( .A(fu_LIFTING_N74), .Y(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n82) );
  XOR2X1 fu_LIFTING_U213 ( .A(fu_LIFTING_N672), .B(fu_LIFTING_N673), .Y(
        fu_LIFTING_n91) );
  NAND2X2 fu_LIFTING_U212 ( .A(fu_LIFTING_n390), .B(fu_LIFTING_n389), .Y(
        fu_LIFTING_n486) );
  INVX2 fu_LIFTING_U211 ( .A(fu_LIFTING_N672), .Y(fu_LIFTING_n262) );
  INVX2 fu_LIFTING_U210 ( .A(fu_LIFTING_N673), .Y(fu_LIFTING_n266) );
  AOI222X2 fu_LIFTING_U209 ( .A0(fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_6_), 
        .A1(fu_LIFTING_n75), .B0(fu_LIFTING_n243), .B1(
        fu_LIFTING_reg_out_tmp_6_), .C0(fu_LIFTING_n246), .C1(
        ic_socket_LIFTING_o1_data0_wire[6]), .Y(fu_LIFTING_n417) );
  AOI222X2 fu_LIFTING_U208 ( .A0(fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_7_), 
        .A1(fu_LIFTING_n242), .B0(fu_LIFTING_n243), .B1(
        fu_LIFTING_reg_out_tmp_7_), .C0(fu_LIFTING_n246), .C1(
        ic_socket_LIFTING_o1_data0_wire[7]), .Y(fu_LIFTING_n418) );
  NAND2X2 fu_LIFTING_U207 ( .A(fu_LIFTING_n388), .B(fu_LIFTING_n387), .Y(
        fu_LIFTING_n487) );
  NAND2X2 fu_LIFTING_U206 ( .A(fu_LIFTING_n386), .B(fu_LIFTING_n385), .Y(
        fu_LIFTING_n488) );
  AOI222X2 fu_LIFTING_U205 ( .A0(fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_8_), 
        .A1(fu_LIFTING_n242), .B0(fu_LIFTING_n243), .B1(
        fu_LIFTING_reg_out_tmp_8_), .C0(fu_LIFTING_n246), .C1(
        ic_socket_LIFTING_o1_data0_wire[8]), .Y(fu_LIFTING_n419) );
  AOI222X2 fu_LIFTING_U204 ( .A0(fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_9_), 
        .A1(fu_LIFTING_n242), .B0(fu_LIFTING_n243), .B1(
        fu_LIFTING_reg_out_tmp_9_), .C0(fu_LIFTING_n246), .C1(
        ic_socket_LIFTING_o1_data0_wire[9]), .Y(fu_LIFTING_n420) );
  ADDFX2 fu_LIFTING_U203 ( .A(fu_LIFTING_mult_79_DP_OP_279_6650_2_n34), .B(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n35), .CI(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n5), .CO(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n4), .S(fu_LIFTING_N188) );
  OAI211X2 fu_LIFTING_U202 ( .A0(fu_LIFTING_n262), .A1(fu_LIFTING_n1), .B0(
        fu_LIFTING_n261), .C0(fu_LIFTING_n260), .Y(fu_LIFTING_n474) );
  AOI222X2 fu_LIFTING_U201 ( .A0(fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_10_), 
        .A1(fu_LIFTING_n242), .B0(fu_LIFTING_n243), .B1(
        fu_LIFTING_reg_out_tmp_10_), .C0(fu_LIFTING_n246), .C1(
        ic_socket_LIFTING_o1_data0_wire[10]), .Y(fu_LIFTING_n421) );
  AOI222X2 fu_LIFTING_U200 ( .A0(fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_11_), 
        .A1(fu_LIFTING_n242), .B0(fu_LIFTING_n74), .B1(
        fu_LIFTING_reg_out_tmp_11_), .C0(fu_LIFTING_n246), .C1(
        ic_socket_LIFTING_o1_data0_wire[11]), .Y(fu_LIFTING_n422) );
  ADDFX2 fu_LIFTING_U199 ( .A(fu_LIFTING_mult_92_DP_OP_280_6650_5_n40), .B(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n41), .CI(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n6), .CO(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n5), .S(fu_LIFTING_N547) );
  ADDFX2 fu_LIFTING_U198 ( .A(fu_LIFTING_mult_79_DP_OP_279_6650_2_n30), .B(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n31), .CI(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n3), .CO(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n2), .S(fu_LIFTING_N190) );
  ADDFX2 fu_LIFTING_U197 ( .A(fu_LIFTING_mult_92_DP_OP_280_6650_5_n38), .B(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n39), .CI(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n5), .CO(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n4), .S(fu_LIFTING_N548) );
  ADDFX2 fu_LIFTING_U196 ( .A(fu_LIFTING_mult_88_DP_OP_277_6650_4_n33), .B(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n34), .CI(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n4), .CO(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n3), .S(fu_LIFTING_N429) );
  ADDFX4 fu_LIFTING_U195 ( .A(fu_LIFTING_mult_96_DP_OP_281_6650_6_n40), .B(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n41), .CI(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n6), .CO(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n5), .S(fu_LIFTING_N667) );
  ADDFX4 fu_LIFTING_U194 ( .A(fu_LIFTING_mult_84_DP_OP_276_6650_3_n32), .B(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n33), .CI(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n3), .CO(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n2), .S(fu_LIFTING_N310) );
  XOR3X4 fu_LIFTING_U193 ( .A(fu_LIFTING_mult_84_DP_OP_276_6650_3_n31), .B(
        fu_LIFTING_n109), .C(fu_LIFTING_n108), .Y(fu_LIFTING_N311) );
  XOR3X4 fu_LIFTING_U192 ( .A(fu_LIFTING_n91), .B(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n2), .C(fu_LIFTING_n90), .Y(
        fu_LIFTING_n92) );
  XOR2X4 fu_LIFTING_U191 ( .A(fu_LIFTING_n93), .B(fu_LIFTING_n92), .Y(
        fu_LIFTING_N71) );
  ADDFX4 fu_LIFTING_U190 ( .A(fu_LIFTING_sub_98_DP_OP_282_1544_7_n45), .B(
        fu_LIFTING_n468), .CI(fu_LIFTING_sub_98_DP_OP_282_1544_7_n8), .CO(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n7), .S(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_25_) );
  CLKBUFX32 fu_LIFTING_U189 ( .A(fu_LIFTING_in2_load_wire), .Y(fu_LIFTING_n248) );
  INVX16 fu_LIFTING_U188 ( .A(n1757), .Y(fu_LIFTING_n42) );
  NOR2X5 fu_LIFTING_U187 ( .A(fu_LIFTING_n72), .B(n1757), .Y(fu_LIFTING_N961)
         );
  ADDFX1 fu_LIFTING_U186 ( .A(fu_LIFTING_N645), .B(fu_LIFTING_N97), .CI(
        fu_LIFTING_N644), .CO(fu_LIFTING_mult_88_DP_OP_277_6650_4_n76), .S(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n77) );
  ADDFX2 fu_LIFTING_U185 ( .A(fu_LIFTING_N702), .B(fu_LIFTING_N698), .CI(
        fu_LIFTING_N701), .CO(fu_LIFTING_mult_84_DP_OP_276_6650_3_n81), .S(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n82) );
  ADDFX2 fu_LIFTING_U184 ( .A(fu_LIFTING_N701), .B(fu_LIFTING_N697), .CI(
        fu_LIFTING_N700), .CO(fu_LIFTING_mult_84_DP_OP_276_6650_3_n79), .S(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n80) );
  ADDFX1 fu_LIFTING_U183 ( .A(fu_LIFTING_N644), .B(fu_LIFTING_N95), .CI(
        fu_LIFTING_N99), .CO(fu_LIFTING_mult_79_DP_OP_279_6650_2_n71), .S(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n72) );
  ADDFX1 fu_LIFTING_U182 ( .A(fu_LIFTING_N99), .B(fu_LIFTING_N95), .CI(
        fu_LIFTING_N98), .CO(fu_LIFTING_mult_88_DP_OP_277_6650_4_n72), .S(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n73) );
  ADDFX1 fu_LIFTING_U181 ( .A(fu_LIFTING_N645), .B(fu_LIFTING_N96), .CI(
        fu_LIFTING_N644), .CO(fu_LIFTING_mult_79_DP_OP_279_6650_2_n73), .S(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n74) );
  ADDFX1 fu_LIFTING_U180 ( .A(fu_LIFTING_N644), .B(fu_LIFTING_N96), .CI(
        fu_LIFTING_N99), .CO(fu_LIFTING_mult_88_DP_OP_277_6650_4_n74), .S(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n75) );
  ADDFX1 fu_LIFTING_U179 ( .A(fu_LIFTING_N98), .B(fu_LIFTING_N94), .CI(
        fu_LIFTING_N97), .CO(fu_LIFTING_mult_88_DP_OP_277_6650_4_n70), .S(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n71) );
  OAI211X2 fu_LIFTING_U178 ( .A0(fu_LIFTING_n76), .A1(fu_LIFTING_n241), .B0(
        fu_LIFTING_n357), .C0(fu_LIFTING_n356), .Y(fu_LIFTING_n444) );
  OAI211X2 fu_LIFTING_U177 ( .A0(fu_LIFTING_n80), .A1(fu_LIFTING_n241), .B0(
        fu_LIFTING_n338), .C0(fu_LIFTING_n337), .Y(fu_LIFTING_n449) );
  OAI211X2 fu_LIFTING_U176 ( .A0(fu_LIFTING_n81), .A1(fu_LIFTING_n1), .B0(
        fu_LIFTING_n332), .C0(fu_LIFTING_n331), .Y(fu_LIFTING_n451) );
  OAI211X2 fu_LIFTING_U175 ( .A0(fu_LIFTING_n78), .A1(fu_LIFTING_n236), .B0(
        fu_LIFTING_n346), .C0(fu_LIFTING_n345), .Y(fu_LIFTING_n447) );
  OAI211X2 fu_LIFTING_U174 ( .A0(fu_LIFTING_n73), .A1(fu_LIFTING_n241), .B0(
        fu_LIFTING_n342), .C0(fu_LIFTING_n341), .Y(fu_LIFTING_n448) );
  ADDFX1 fu_LIFTING_U173 ( .A(fu_LIFTING_N99), .B(fu_LIFTING_n69), .CI(
        fu_LIFTING_N96), .CO(fu_LIFTING_mult_96_DP_OP_281_6650_6_n71), .S(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n72) );
  NAND2X2 fu_LIFTING_U172 ( .A(fu_LIFTING_n77), .B(fu_LIFTING_n3), .Y(
        fu_LIFTING_n88) );
  OAI211X2 fu_LIFTING_U171 ( .A0(fu_LIFTING_n82), .A1(fu_LIFTING_n2), .B0(
        fu_LIFTING_n335), .C0(fu_LIFTING_n334), .Y(fu_LIFTING_n450) );
  OAI211X2 fu_LIFTING_U170 ( .A0(fu_LIFTING_n71), .A1(fu_LIFTING_n1), .B0(
        fu_LIFTING_n329), .C0(fu_LIFTING_n328), .Y(fu_LIFTING_n452) );
  ADDFX1 fu_LIFTING_U169 ( .A(fu_LIFTING_N96), .B(fu_LIFTING_N91), .CI(
        fu_LIFTING_N95), .CO(fu_LIFTING_mult_79_DP_OP_279_6650_2_n63), .S(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n64) );
  NAND2X2 fu_LIFTING_U168 ( .A(fu_LIFTING_n77), .B(fu_LIFTING_N647), .Y(
        fu_LIFTING_n89) );
  OAI211X2 fu_LIFTING_U167 ( .A0(fu_LIFTING_n68), .A1(fu_LIFTING_n241), .B0(
        fu_LIFTING_n326), .C0(fu_LIFTING_n325), .Y(fu_LIFTING_n453) );
  OAI21X4 fu_LIFTING_U166 ( .A0(fu_LIFTING_N703), .A1(fu_LIFTING_n127), .B0(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n82), .Y(fu_LIFTING_n126) );
  ADDFX1 fu_LIFTING_U165 ( .A(fu_LIFTING_N95), .B(fu_LIFTING_N90), .CI(
        fu_LIFTING_N94), .CO(fu_LIFTING_mult_79_DP_OP_279_6650_2_n61), .S(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n62) );
  OAI21X4 fu_LIFTING_U164 ( .A0(fu_LIFTING_mult_88_DP_OP_277_6650_4_n78), .A1(
        fu_LIFTING_n121), .B0(fu_LIFTING_mult_88_DP_OP_277_6650_4_n77), .Y(
        fu_LIFTING_n120) );
  OAI21X4 fu_LIFTING_U163 ( .A0(fu_LIFTING_mult_84_DP_OP_276_6650_3_n81), .A1(
        fu_LIFTING_n113), .B0(fu_LIFTING_mult_84_DP_OP_276_6650_3_n80), .Y(
        fu_LIFTING_n112) );
  OAI211X2 fu_LIFTING_U162 ( .A0(fu_LIFTING_n67), .A1(fu_LIFTING_n1), .B0(
        fu_LIFTING_n323), .C0(fu_LIFTING_n322), .Y(fu_LIFTING_n454) );
  OAI211X2 fu_LIFTING_U161 ( .A0(fu_LIFTING_n70), .A1(fu_LIFTING_n2), .B0(
        fu_LIFTING_n360), .C0(fu_LIFTING_n359), .Y(fu_LIFTING_n443) );
  ADDFX1 fu_LIFTING_U160 ( .A(fu_LIFTING_N92), .B(fu_LIFTING_N87), .CI(
        fu_LIFTING_N91), .CO(fu_LIFTING_mult_79_DP_OP_279_6650_2_n55), .S(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n56) );
  OAI211X2 fu_LIFTING_U159 ( .A0(fu_LIFTING_n66), .A1(fu_LIFTING_n1), .B0(
        fu_LIFTING_n320), .C0(fu_LIFTING_n319), .Y(fu_LIFTING_n455) );
  OAI211X2 fu_LIFTING_U158 ( .A0(fu_LIFTING_n65), .A1(fu_LIFTING_n236), .B0(
        fu_LIFTING_n317), .C0(fu_LIFTING_n316), .Y(fu_LIFTING_n456) );
  OAI21X4 fu_LIFTING_U157 ( .A0(fu_LIFTING_mult_75_DP_OP_278_6650_1_n111), 
        .A1(fu_LIFTING_n100), .B0(fu_LIFTING_mult_75_DP_OP_278_6650_1_n110), 
        .Y(fu_LIFTING_n99) );
  ADDFX1 fu_LIFTING_U156 ( .A(fu_LIFTING_N89), .B(fu_LIFTING_N85), .CI(
        fu_LIFTING_N88), .CO(fu_LIFTING_mult_88_DP_OP_277_6650_4_n52), .S(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n53) );
  OAI211X2 fu_LIFTING_U155 ( .A0(fu_LIFTING_n61), .A1(fu_LIFTING_n1), .B0(
        fu_LIFTING_n314), .C0(fu_LIFTING_n313), .Y(fu_LIFTING_n457) );
  OAI211X2 fu_LIFTING_U154 ( .A0(fu_LIFTING_n63), .A1(fu_LIFTING_n241), .B0(
        fu_LIFTING_n311), .C0(fu_LIFTING_n310), .Y(fu_LIFTING_n458) );
  ADDFX1 fu_LIFTING_U153 ( .A(fu_LIFTING_N90), .B(fu_LIFTING_N85), .CI(
        fu_LIFTING_N89), .CO(fu_LIFTING_mult_79_DP_OP_279_6650_2_n51), .S(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n52) );
  OAI211X2 fu_LIFTING_U152 ( .A0(fu_LIFTING_n60), .A1(fu_LIFTING_n1), .B0(
        fu_LIFTING_n308), .C0(fu_LIFTING_n307), .Y(fu_LIFTING_n459) );
  OAI211X2 fu_LIFTING_U151 ( .A0(fu_LIFTING_n59), .A1(fu_LIFTING_n1), .B0(
        fu_LIFTING_n305), .C0(fu_LIFTING_n304), .Y(fu_LIFTING_n460) );
  ADDFX1 fu_LIFTING_U150 ( .A(fu_LIFTING_N687), .B(fu_LIFTING_N683), .CI(
        fu_LIFTING_N686), .CO(fu_LIFTING_mult_84_DP_OP_276_6650_3_n51), .S(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n52) );
  OAI211X2 fu_LIFTING_U149 ( .A0(fu_LIFTING_n58), .A1(fu_LIFTING_n236), .B0(
        fu_LIFTING_n302), .C0(fu_LIFTING_n301), .Y(fu_LIFTING_n461) );
  OAI211X2 fu_LIFTING_U148 ( .A0(fu_LIFTING_n56), .A1(fu_LIFTING_n1), .B0(
        fu_LIFTING_n299), .C0(fu_LIFTING_n298), .Y(fu_LIFTING_n462) );
  ADDFX4 fu_LIFTING_U147 ( .A(fu_LIFTING_mult_75_DP_OP_278_6650_1_n98), .B(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n100), .CI(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n23), .CO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n22), .S(fu_LIFTING_N50) );
  OAI211X2 fu_LIFTING_U146 ( .A0(fu_LIFTING_n55), .A1(fu_LIFTING_n1), .B0(
        fu_LIFTING_n296), .C0(fu_LIFTING_n295), .Y(fu_LIFTING_n463) );
  INVX4 fu_LIFTING_U145 ( .A(fu_LIFTING_N680), .Y(fu_LIFTING_n52) );
  INVX2 fu_LIFTING_U144 ( .A(fu_LIFTING_N80), .Y(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n88) );
  ADDFHX2 fu_LIFTING_U143 ( .A(fu_LIFTING_mult_75_DP_OP_278_6650_1_n95), .B(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n22), .CI(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n97), .CO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n21), .S(fu_LIFTING_N51) );
  ADDFX2 fu_LIFTING_U142 ( .A(fu_LIFTING_mult_96_DP_OP_281_6650_6_n70), .B(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n71), .CI(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n21), .CO(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n20), .S(fu_LIFTING_N652) );
  OAI211X2 fu_LIFTING_U141 ( .A0(fu_LIFTING_n54), .A1(fu_LIFTING_n1), .B0(
        fu_LIFTING_n293), .C0(fu_LIFTING_n292), .Y(fu_LIFTING_n464) );
  INVX4 fu_LIFTING_U140 ( .A(fu_LIFTING_N678), .Y(fu_LIFTING_n49) );
  OAI211X2 fu_LIFTING_U139 ( .A0(fu_LIFTING_n53), .A1(fu_LIFTING_n1), .B0(
        fu_LIFTING_n290), .C0(fu_LIFTING_n289), .Y(fu_LIFTING_n465) );
  ADDFX1 fu_LIFTING_U138 ( .A(fu_LIFTING_N84), .B(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n86), .CI(fu_LIFTING_N81), .CO(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n41), .S(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n42) );
  ADDFX1 fu_LIFTING_U137 ( .A(fu_LIFTING_N81), .B(fu_LIFTING_N77), .CI(
        fu_LIFTING_N80), .CO(fu_LIFTING_mult_88_DP_OP_277_6650_4_n36), .S(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n37) );
  CLKXOR2X2 fu_LIFTING_U136 ( .A(fu_LIFTING_n41), .B(fu_LIFTING_n479), .Y(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n68) );
  ADDFX1 fu_LIFTING_U135 ( .A(fu_LIFTING_N83), .B(fu_LIFTING_n48), .CI(
        fu_LIFTING_N80), .CO(fu_LIFTING_mult_96_DP_OP_281_6650_6_n39), .S(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n40) );
  OAI211X2 fu_LIFTING_U134 ( .A0(fu_LIFTING_n51), .A1(fu_LIFTING_n236), .B0(
        fu_LIFTING_n284), .C0(fu_LIFTING_n283), .Y(fu_LIFTING_n467) );
  CLKXOR2X2 fu_LIFTING_U133 ( .A(fu_LIFTING_n41), .B(fu_LIFTING_n480), .Y(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n67) );
  ADDFX1 fu_LIFTING_U132 ( .A(fu_LIFTING_N81), .B(fu_LIFTING_N76), .CI(
        fu_LIFTING_N80), .CO(fu_LIFTING_mult_79_DP_OP_279_6650_2_n33), .S(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n34) );
  ADDFX1 fu_LIFTING_U131 ( .A(fu_LIFTING_N80), .B(fu_LIFTING_N76), .CI(
        fu_LIFTING_N79), .CO(fu_LIFTING_mult_88_DP_OP_277_6650_4_n34), .S(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n35) );
  MX2X4 fu_LIFTING_U130 ( .A(fu_LIFTING_reg_x2_28_), .B(rf_RF_t1data_wire[28]), 
        .S0(fu_LIFTING_n248), .Y(fu_LIFTING_N675) );
  INVX4 fu_LIFTING_U129 ( .A(fu_LIFTING_N676), .Y(fu_LIFTING_n46) );
  AOI22X2 fu_LIFTING_U128 ( .A0(fu_LIFTING_N678), .A1(fu_LIFTING_n46), .B0(
        fu_LIFTING_N676), .B1(fu_LIFTING_n49), .Y(fu_LIFTING_n123) );
  AOI22X2 fu_LIFTING_U127 ( .A0(fu_LIFTING_N79), .A1(fu_LIFTING_n45), .B0(
        fu_LIFTING_N76), .B1(fu_LIFTING_n51), .Y(fu_LIFTING_n131) );
  OAI211X2 fu_LIFTING_U126 ( .A0(fu_LIFTING_n47), .A1(fu_LIFTING_n241), .B0(
        fu_LIFTING_n278), .C0(fu_LIFTING_n277), .Y(fu_LIFTING_n469) );
  MX2X4 fu_LIFTING_U125 ( .A(fu_LIFTING_reg_x2_29_), .B(n1861), .S0(
        fu_LIFTING_n248), .Y(fu_LIFTING_N674) );
  OAI211X2 fu_LIFTING_U124 ( .A0(fu_LIFTING_n46), .A1(fu_LIFTING_n241), .B0(
        fu_LIFTING_n275), .C0(fu_LIFTING_n274), .Y(fu_LIFTING_n470) );
  XNOR2X1 fu_LIFTING_U123 ( .A(fu_LIFTING_mult_75_DP_OP_278_6650_1_n37), .B(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n36), .Y(fu_LIFTING_n93) );
  NAND2X2 fu_LIFTING_U122 ( .A(fu_LIFTING_n382), .B(fu_LIFTING_n381), .Y(
        fu_LIFTING_n490) );
  ADDFX2 fu_LIFTING_U121 ( .A(fu_LIFTING_mult_79_DP_OP_279_6650_2_n32), .B(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n33), .CI(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n4), .CO(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n3), .S(fu_LIFTING_N189) );
  ADDFX2 fu_LIFTING_U120 ( .A(fu_LIFTING_mult_84_DP_OP_276_6650_3_n40), .B(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n41), .CI(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n7), .CO(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n6), .S(fu_LIFTING_N306) );
  ADDFX2 fu_LIFTING_U119 ( .A(fu_LIFTING_mult_88_DP_OP_277_6650_4_n35), .B(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n36), .CI(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n5), .CO(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n4), .S(fu_LIFTING_N428) );
  ADDFX4 fu_LIFTING_U118 ( .A(fu_LIFTING_mult_84_DP_OP_276_6650_3_n38), .B(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n39), .CI(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n6), .CO(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n5), .S(fu_LIFTING_N307) );
  INVX8 fu_LIFTING_U117 ( .A(fu_LIFTING_n408), .Y(fu_LIFTING_n236) );
  CLKBUFX32 fu_LIFTING_U116 ( .A(fu_LIFTING_sub_98_DP_OP_282_1544_7_n71), .Y(
        fu_LIFTING_n41) );
  MX2X8 fu_LIFTING_U115 ( .A(fu_LIFTING_reg_x1_2_), .B(n1810), .S0(
        fu_LIFTING_n42), .Y(fu_LIFTING_N645) );
  ADDFX1 fu_LIFTING_U114 ( .A(fu_LIFTING_N646), .B(fu_LIFTING_N97), .CI(
        fu_LIFTING_N645), .CO(fu_LIFTING_mult_79_DP_OP_279_6650_2_n75), .S(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n76) );
  ADDFX1 fu_LIFTING_U113 ( .A(fu_LIFTING_N699), .B(fu_LIFTING_n71), .CI(
        fu_LIFTING_N697), .CO(fu_LIFTING_mult_92_DP_OP_280_6650_5_n73), .S(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n74) );
  ADDFX1 fu_LIFTING_U112 ( .A(fu_LIFTING_N698), .B(fu_LIFTING_n68), .CI(
        fu_LIFTING_N696), .CO(fu_LIFTING_mult_92_DP_OP_280_6650_5_n71), .S(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n72) );
  ADDFX1 fu_LIFTING_U111 ( .A(fu_LIFTING_N98), .B(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n100), .CI(fu_LIFTING_N95), .CO(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n69), .S(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n70) );
  ADDFX1 fu_LIFTING_U110 ( .A(fu_LIFTING_N94), .B(fu_LIFTING_n62), .CI(
        fu_LIFTING_N91), .CO(fu_LIFTING_mult_96_DP_OP_281_6650_6_n61), .S(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n62) );
  ADDFX1 fu_LIFTING_U109 ( .A(fu_LIFTING_N93), .B(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n95), .CI(fu_LIFTING_N90), .CO(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n59), .S(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n60) );
  ADDFX2 fu_LIFTING_U108 ( .A(fu_LIFTING_mult_88_DP_OP_277_6650_4_n71), .B(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n72), .CI(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n23), .CO(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n22), .S(fu_LIFTING_N410) );
  ADDFX1 fu_LIFTING_U107 ( .A(fu_LIFTING_N690), .B(fu_LIFTING_n57), .CI(
        fu_LIFTING_N688), .CO(fu_LIFTING_mult_92_DP_OP_280_6650_5_n55), .S(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n56) );
  ADDFX2 fu_LIFTING_U106 ( .A(fu_LIFTING_mult_88_DP_OP_277_6650_4_n69), .B(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n70), .CI(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n22), .CO(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n21), .S(fu_LIFTING_N411) );
  ADDFX1 fu_LIFTING_U105 ( .A(fu_LIFTING_mult_79_DP_OP_279_6650_2_n64), .B(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n65), .CI(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n20), .CO(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n19), .S(fu_LIFTING_N173) );
  ADDFX1 fu_LIFTING_U104 ( .A(fu_LIFTING_N689), .B(fu_LIFTING_n56), .CI(
        fu_LIFTING_N687), .CO(fu_LIFTING_mult_92_DP_OP_280_6650_5_n53), .S(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n54) );
  ADDFX2 fu_LIFTING_U103 ( .A(fu_LIFTING_mult_92_DP_OP_280_6650_5_n70), .B(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n71), .CI(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n21), .CO(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n20), .S(fu_LIFTING_N532) );
  ADDFX2 fu_LIFTING_U102 ( .A(fu_LIFTING_mult_79_DP_OP_279_6650_2_n54), .B(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n55), .CI(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n15), .CO(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n14), .S(fu_LIFTING_N178) );
  ADDFX2 fu_LIFTING_U101 ( .A(fu_LIFTING_mult_96_DP_OP_281_6650_6_n68), .B(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n69), .CI(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n20), .CO(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n19), .S(fu_LIFTING_N653) );
  ADDFX1 fu_LIFTING_U100 ( .A(fu_LIFTING_N681), .B(fu_LIFTING_N677), .CI(
        fu_LIFTING_N680), .CO(fu_LIFTING_mult_84_DP_OP_276_6650_3_n39), .S(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n40) );
  ADDFX2 fu_LIFTING_U99 ( .A(fu_LIFTING_mult_79_DP_OP_279_6650_2_n50), .B(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n51), .CI(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n13), .CO(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n12), .S(fu_LIFTING_N180) );
  MX2X4 fu_LIFTING_U98 ( .A(fu_LIFTING_reg_x1_28_), .B(rf_RF_t1data_wire[28]), 
        .S0(fu_LIFTING_n249), .Y(fu_LIFTING_N75) );
  MX2X4 fu_LIFTING_U97 ( .A(fu_LIFTING_reg_x1_29_), .B(n1861), .S0(
        fu_LIFTING_n249), .Y(fu_LIFTING_N74) );
  ADDFX2 fu_LIFTING_U96 ( .A(fu_LIFTING_mult_88_DP_OP_277_6650_4_n51), .B(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n52), .CI(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n13), .CO(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n12), .S(fu_LIFTING_N420) );
  ADDFX2 fu_LIFTING_U95 ( .A(fu_LIFTING_mult_96_DP_OP_281_6650_6_n60), .B(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n61), .CI(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n16), .CO(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n15), .S(fu_LIFTING_N657) );
  ADDFX2 fu_LIFTING_U94 ( .A(fu_LIFTING_mult_96_DP_OP_281_6650_6_n58), .B(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n59), .CI(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n15), .CO(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n14), .S(fu_LIFTING_N658) );
  ADDFX2 fu_LIFTING_U93 ( .A(fu_LIFTING_mult_84_DP_OP_276_6650_3_n50), .B(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n51), .CI(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n12), .CO(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n11), .S(fu_LIFTING_N301) );
  NAND2X2 fu_LIFTING_U92 ( .A(fu_LIFTING_n380), .B(fu_LIFTING_n379), .Y(
        fu_LIFTING_n491) );
  NAND2X2 fu_LIFTING_U91 ( .A(fu_LIFTING_n378), .B(fu_LIFTING_n377), .Y(
        fu_LIFTING_n492) );
  ADDFX2 fu_LIFTING_U90 ( .A(fu_LIFTING_mult_88_DP_OP_277_6650_4_n31), .B(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n32), .CI(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n3), .CO(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n2), .S(fu_LIFTING_N430) );
  NAND2X2 fu_LIFTING_U89 ( .A(fu_LIFTING_n376), .B(fu_LIFTING_n375), .Y(
        fu_LIFTING_n493) );
  ADDFX2 fu_LIFTING_U88 ( .A(fu_LIFTING_mult_92_DP_OP_280_6650_5_n34), .B(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n35), .CI(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n3), .CO(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n2), .S(fu_LIFTING_N550) );
  AOI222X2 fu_LIFTING_U87 ( .A0(fu_LIFTING_N668), .A1(fu_LIFTING_n240), .B0(
        fu_LIFTING_n37), .B1(fu_LIFTING_N548), .C0(fu_LIFTING_n238), .C1(
        fu_LIFTING_N188), .Y(fu_LIFTING_n367) );
  XOR3X2 fu_LIFTING_U86 ( .A(fu_LIFTING_mult_88_DP_OP_277_6650_4_n30), .B(
        fu_LIFTING_n117), .C(fu_LIFTING_n116), .Y(fu_LIFTING_N431) );
  AOI222X2 fu_LIFTING_U85 ( .A0(fu_LIFTING_N67), .A1(fu_LIFTING_n36), .B0(
        fu_LIFTING_n83), .B1(fu_LIFTING_N427), .C0(fu_LIFTING_n235), .C1(
        fu_LIFTING_N307), .Y(fu_LIFTING_n370) );
  AOI222X2 fu_LIFTING_U84 ( .A0(fu_LIFTING_N669), .A1(fu_LIFTING_n240), .B0(
        fu_LIFTING_n37), .B1(fu_LIFTING_N549), .C0(fu_LIFTING_n238), .C1(
        fu_LIFTING_N189), .Y(fu_LIFTING_n365) );
  AOI222X2 fu_LIFTING_U83 ( .A0(fu_LIFTING_N68), .A1(fu_LIFTING_n36), .B0(
        fu_LIFTING_n83), .B1(fu_LIFTING_N428), .C0(fu_LIFTING_n235), .C1(
        fu_LIFTING_N308), .Y(fu_LIFTING_n368) );
  XOR3X2 fu_LIFTING_U82 ( .A(fu_LIFTING_n123), .B(fu_LIFTING_n122), .C(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n33), .Y(fu_LIFTING_N551) );
  AOI222X2 fu_LIFTING_U81 ( .A0(fu_LIFTING_N670), .A1(fu_LIFTING_n240), .B0(
        fu_LIFTING_n234), .B1(fu_LIFTING_N310), .C0(fu_LIFTING_n238), .C1(
        fu_LIFTING_N190), .Y(fu_LIFTING_n363) );
  AOI222X2 fu_LIFTING_U80 ( .A0(fu_LIFTING_N70), .A1(fu_LIFTING_n36), .B0(
        fu_LIFTING_n83), .B1(fu_LIFTING_N430), .C0(fu_LIFTING_n37), .C1(
        fu_LIFTING_N550), .Y(fu_LIFTING_n364) );
  CLKBUFX6 fu_LIFTING_U79 ( .A(n2211), .Y(fu_LIFTING_n247) );
  CLKINVX32 fu_LIFTING_U78 ( .A(fu_LIFTING_n2), .Y(fu_LIFTING_n83) );
  CLKMX2X8 fu_LIFTING_U77 ( .A(fu_LIFTING_reg_x2_8_), .B(rf_RF_t1data_wire[8]), 
        .S0(fu_LIFTING_n248), .Y(fu_LIFTING_N695) );
  CLKMX2X8 fu_LIFTING_U75 ( .A(fu_LIFTING_reg_x1_6_), .B(n1818), .S0(
        fu_LIFTING_n42), .Y(fu_LIFTING_N97) );
  CLKMX2X8 fu_LIFTING_U74 ( .A(fu_LIFTING_reg_x2_7_), .B(n1814), .S0(
        fu_LIFTING_n248), .Y(fu_LIFTING_N696) );
  INVX4 fu_LIFTING_U73 ( .A(fu_LIFTING_N645), .Y(fu_LIFTING_n39) );
  CLKMX2X8 fu_LIFTING_U72 ( .A(fu_LIFTING_reg_x2_11_), .B(
        rf_RF_t1data_wire[11]), .S0(fu_LIFTING_n248), .Y(fu_LIFTING_N692) );
  CLKMX2X8 fu_LIFTING_U71 ( .A(fu_LIFTING_reg_x2_12_), .B(n1820), .S0(
        fu_LIFTING_n248), .Y(fu_LIFTING_N691) );
  INVX4 fu_LIFTING_U70 ( .A(fu_LIFTING_N703), .Y(fu_LIFTING_n70) );
  INVX2 fu_LIFTING_U69 ( .A(fu_LIFTING_N90), .Y(fu_LIFTING_n65) );
  INVX2 fu_LIFTING_U68 ( .A(fu_LIFTING_N690), .Y(fu_LIFTING_n64) );
  CLKMX2X8 fu_LIFTING_U67 ( .A(fu_LIFTING_reg_x2_14_), .B(
        rf_RF_t1data_wire[14]), .S0(fu_LIFTING_n248), .Y(fu_LIFTING_N689) );
  CLKMX2X8 fu_LIFTING_U66 ( .A(fu_LIFTING_reg_x2_16_), .B(
        rf_RF_t1data_wire[16]), .S0(fu_LIFTING_n248), .Y(fu_LIFTING_N687) );
  INVX2 fu_LIFTING_U65 ( .A(fu_LIFTING_N88), .Y(fu_LIFTING_n62) );
  CLKMX2X8 fu_LIFTING_U64 ( .A(fu_LIFTING_reg_x2_17_), .B(
        rf_RF_t1data_wire[17]), .S0(fu_LIFTING_n248), .Y(fu_LIFTING_N686) );
  INVX2 fu_LIFTING_U63 ( .A(fu_LIFTING_N685), .Y(fu_LIFTING_n57) );
  CLKMX2X8 fu_LIFTING_U62 ( .A(fu_LIFTING_reg_x2_19_), .B(
        rf_RF_t1data_wire[19]), .S0(fu_LIFTING_n248), .Y(fu_LIFTING_N684) );
  INVX2 fu_LIFTING_U61 ( .A(fu_LIFTING_N85), .Y(fu_LIFTING_n58) );
  CLKMX2X8 fu_LIFTING_U60 ( .A(fu_LIFTING_reg_x2_20_), .B(
        rf_RF_t1data_wire[20]), .S0(fu_LIFTING_n248), .Y(fu_LIFTING_N683) );
  CLKMX2X8 fu_LIFTING_U59 ( .A(fu_LIFTING_reg_x2_21_), .B(
        rf_RF_t1data_wire[21]), .S0(fu_LIFTING_n248), .Y(fu_LIFTING_N682) );
  CLKMX2X8 fu_LIFTING_U58 ( .A(fu_LIFTING_reg_x2_22_), .B(
        rf_RF_t1data_wire[22]), .S0(fu_LIFTING_n248), .Y(fu_LIFTING_N681) );
  AOI222X2 fu_LIFTING_U57 ( .A0(fu_LIFTING_N48), .A1(fu_LIFTING_n36), .B0(
        fu_LIFTING_n234), .B1(fu_LIFTING_N288), .C0(fu_LIFTING_n238), .C1(
        fu_LIFTING_N168), .Y(fu_LIFTING_n410) );
  CLKMX2X8 fu_LIFTING_U56 ( .A(fu_LIFTING_reg_x2_23_), .B(
        rf_RF_t1data_wire[23]), .S0(fu_LIFTING_n248), .Y(fu_LIFTING_N680) );
  AOI222X2 fu_LIFTING_U55 ( .A0(fu_LIFTING_N650), .A1(fu_LIFTING_n240), .B0(
        fu_LIFTING_n234), .B1(fu_LIFTING_N290), .C0(fu_LIFTING_n238), .C1(
        fu_LIFTING_N170), .Y(fu_LIFTING_n403) );
  CLKMX2X8 fu_LIFTING_U54 ( .A(fu_LIFTING_reg_x1_25_), .B(
        rf_RF_t1data_wire[25]), .S0(fu_LIFTING_n249), .Y(fu_LIFTING_N78) );
  INVX2 fu_LIFTING_U53 ( .A(fu_LIFTING_N679), .Y(fu_LIFTING_n50) );
  CLKMX2X8 fu_LIFTING_U52 ( .A(fu_LIFTING_reg_x1_26_), .B(
        rf_RF_t1data_wire[26]), .S0(fu_LIFTING_n249), .Y(fu_LIFTING_N77) );
  CLKMX2X8 fu_LIFTING_U51 ( .A(fu_LIFTING_reg_x2_26_), .B(
        rf_RF_t1data_wire[26]), .S0(fu_LIFTING_n248), .Y(fu_LIFTING_N677) );
  CLKMX2X8 fu_LIFTING_U50 ( .A(fu_LIFTING_reg_x2_27_), .B(
        rf_RF_t1data_wire[27]), .S0(fu_LIFTING_n248), .Y(fu_LIFTING_N676) );
  CLKMX2X6 fu_LIFTING_U49 ( .A(fu_LIFTING_reg_x1_27_), .B(
        rf_RF_t1data_wire[27]), .S0(fu_LIFTING_n249), .Y(fu_LIFTING_N76) );
  ADDFX2 fu_LIFTING_U48 ( .A(fu_LIFTING_mult_92_DP_OP_280_6650_5_n54), .B(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n55), .CI(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n13), .CO(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n12), .S(fu_LIFTING_N540) );
  ADDFX2 fu_LIFTING_U47 ( .A(fu_LIFTING_mult_92_DP_OP_280_6650_5_n52), .B(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n53), .CI(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n12), .CO(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n11), .S(fu_LIFTING_N541) );
  XNOR2X2 fu_LIFTING_U46 ( .A(fu_LIFTING_N73), .B(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n2), .Y(fu_LIFTING_n104) );
  NAND2X2 fu_LIFTING_U45 ( .A(fu_LIFTING_n374), .B(fu_LIFTING_n373), .Y(
        fu_LIFTING_n494) );
  NAND2X2 fu_LIFTING_U44 ( .A(fu_LIFTING_n372), .B(fu_LIFTING_n371), .Y(
        fu_LIFTING_n495) );
  AOI222X2 fu_LIFTING_U43 ( .A0(fu_LIFTING_N69), .A1(fu_LIFTING_n36), .B0(
        fu_LIFTING_n83), .B1(fu_LIFTING_N429), .C0(fu_LIFTING_n235), .C1(
        fu_LIFTING_N309), .Y(fu_LIFTING_n366) );
  CLKXOR2X4 fu_LIFTING_U42 ( .A(fu_LIFTING_N73), .B(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n2), .Y(fu_LIFTING_n130) );
  NAND2X2 fu_LIFTING_U41 ( .A(fu_LIFTING_n368), .B(fu_LIFTING_n367), .Y(
        fu_LIFTING_n497) );
  NAND2X2 fu_LIFTING_U40 ( .A(fu_LIFTING_n366), .B(fu_LIFTING_n365), .Y(
        fu_LIFTING_n498) );
  NAND2X2 fu_LIFTING_U39 ( .A(fu_LIFTING_n364), .B(fu_LIFTING_n363), .Y(
        fu_LIFTING_n499) );
  AOI222X2 fu_LIFTING_U38 ( .A0(fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_29_), 
        .A1(fu_LIFTING_n242), .B0(fu_LIFTING_n243), .B1(
        fu_LIFTING_reg_out_tmp_29_), .C0(fu_LIFTING_n246), .C1(
        ic_socket_LIFTING_o1_data0_wire[29]), .Y(fu_LIFTING_n440) );
  CLKINVX40 fu_LIFTING_U37 ( .A(fu_LIFTING_n237), .Y(fu_LIFTING_n37) );
  CLKINVX40 fu_LIFTING_U36 ( .A(fu_LIFTING_n236), .Y(fu_LIFTING_n36) );
  CLKMX2X8 fu_LIFTING_U35 ( .A(fu_LIFTING_reg_x1_3_), .B(rf_RF_t1data_wire[3]), 
        .S0(fu_LIFTING_n42), .Y(fu_LIFTING_N644) );
  CLKMX2X8 fu_LIFTING_U34 ( .A(fu_LIFTING_reg_x2_9_), .B(n1812), .S0(
        fu_LIFTING_n248), .Y(fu_LIFTING_N694) );
  CLKMX2X8 fu_LIFTING_U33 ( .A(fu_LIFTING_reg_x2_25_), .B(
        rf_RF_t1data_wire[25]), .S0(fu_LIFTING_n248), .Y(fu_LIFTING_N678) );
  ADDHX2 fu_LIFTING_U32 ( .A(fu_LIFTING_n79), .B(fu_LIFTING_N644), .CO(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n79), .S(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n80) );
  AND2X2 fu_LIFTING_U31 ( .A(fu_LIFTING_n40), .B(fu_LIFTING_n39), .Y(
        fu_LIFTING_n3) );
  CLKMX2X6 fu_LIFTING_U30 ( .A(fu_LIFTING_reg_x1_0_), .B(n2111), .S0(
        fu_LIFTING_n42), .Y(fu_LIFTING_N647) );
  OAI21X4 fu_LIFTING_U29 ( .A0(fu_LIFTING_n87), .A1(fu_LIFTING_n102), .B0(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n107), .Y(fu_LIFTING_n101) );
  CLKXOR2X4 fu_LIFTING_U28 ( .A(fu_LIFTING_n41), .B(fu_LIFTING_n500), .Y(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n46) );
  ADDFHX2 fu_LIFTING_U27 ( .A(fu_LIFTING_mult_75_DP_OP_278_6650_1_n101), .B(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n103), .CI(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n24), .CO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n23), .S(fu_LIFTING_N49) );
  ADDFHX2 fu_LIFTING_U26 ( .A(fu_LIFTING_mult_75_DP_OP_278_6650_1_n59), .B(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n61), .CI(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n10), .CO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n9), .S(fu_LIFTING_N63) );
  CLKXOR2X2 fu_LIFTING_U25 ( .A(fu_LIFTING_n41), .B(fu_LIFTING_n499), .Y(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n48) );
  ADDFX2 fu_LIFTING_U24 ( .A(fu_LIFTING_sub_98_DP_OP_282_1544_7_n48), .B(
        fu_LIFTING_n465), .CI(fu_LIFTING_sub_98_DP_OP_282_1544_7_n11), .CO(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n10), .S(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_22_) );
  NAND2X2 fu_LIFTING_U23 ( .A(fu_LIFTING_n370), .B(fu_LIFTING_n369), .Y(
        fu_LIFTING_n496) );
  ADDFX2 fu_LIFTING_U22 ( .A(fu_LIFTING_sub_98_DP_OP_282_1544_7_n51), .B(
        fu_LIFTING_n462), .CI(fu_LIFTING_sub_98_DP_OP_282_1544_7_n14), .CO(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n13), .S(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_19_) );
  CLKXOR2X2 fu_LIFTING_U21 ( .A(fu_LIFTING_n41), .B(fu_LIFTING_n493), .Y(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n54) );
  ADDFX2 fu_LIFTING_U20 ( .A(fu_LIFTING_mult_96_DP_OP_281_6650_6_n34), .B(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n35), .CI(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n3), .CO(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n2), .S(fu_LIFTING_N670) );
  ADDFX1 fu_LIFTING_U19 ( .A(fu_LIFTING_mult_75_DP_OP_278_6650_1_n38), .B(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n40), .CI(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n3), .CO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n2), .S(fu_LIFTING_N70) );
  ADDFX2 fu_LIFTING_U18 ( .A(fu_LIFTING_mult_96_DP_OP_281_6650_6_n38), .B(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n39), .CI(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n5), .CO(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n4), .S(fu_LIFTING_N668) );
  ADDFX1 fu_LIFTING_U17 ( .A(fu_LIFTING_mult_75_DP_OP_278_6650_1_n44), .B(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n46), .CI(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n5), .CO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n4), .S(fu_LIFTING_N68) );
  ADDFX1 fu_LIFTING_U16 ( .A(fu_LIFTING_mult_75_DP_OP_278_6650_1_n47), .B(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n49), .CI(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n6), .CO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n5), .S(fu_LIFTING_N67) );
  ADDFX1 fu_LIFTING_U15 ( .A(fu_LIFTING_mult_75_DP_OP_278_6650_1_n56), .B(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n58), .CI(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n9), .CO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n8), .S(fu_LIFTING_N64) );
  BUFX8 fu_LIFTING_U14 ( .A(fu_LIFTING_n231), .Y(fu_LIFTING_n237) );
  ADDFX1 fu_LIFTING_U13 ( .A(fu_LIFTING_mult_75_DP_OP_278_6650_1_n68), .B(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n70), .CI(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n13), .CO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n12), .S(fu_LIFTING_N60) );
  CLKMX2X8 fu_LIFTING_U12 ( .A(fu_LIFTING_reg_x1_1_), .B(n2110), .S0(
        fu_LIFTING_n42), .Y(fu_LIFTING_N646) );
  INVX2 fu_LIFTING_U11 ( .A(fu_LIFTING_N646), .Y(fu_LIFTING_n40) );
  CMPR42X1 fu_LIFTING_U10 ( .A(fu_LIFTING_N688), .B(fu_LIFTING_N689), .C(
        fu_LIFTING_N685), .D(fu_LIFTING_N684), .ICI(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n72), .S(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n71), .ICO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n69), .CO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n70) );
  CLKXOR2X2 fu_LIFTING_U9 ( .A(fu_LIFTING_n41), .B(fu_LIFTING_n498), .Y(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n49) );
  CLKXOR2X2 fu_LIFTING_U8 ( .A(fu_LIFTING_n41), .B(fu_LIFTING_n495), .Y(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n52) );
  ADDFX2 fu_LIFTING_U7 ( .A(fu_LIFTING_sub_98_DP_OP_282_1544_7_n52), .B(
        fu_LIFTING_n461), .CI(fu_LIFTING_sub_98_DP_OP_282_1544_7_n15), .CO(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n14), .S(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_18_) );
  CLKXOR2X2 fu_LIFTING_U6 ( .A(fu_LIFTING_n41), .B(fu_LIFTING_n497), .Y(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n50) );
  CLKXOR2X2 fu_LIFTING_U5 ( .A(fu_LIFTING_n41), .B(fu_LIFTING_n494), .Y(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n53) );
  OR2X6 fu_LIFTING_U4 ( .A(fu_LIFTING_n259), .B(fu_LIFTING_n250), .Y(
        fu_LIFTING_n2) );
  INVX20 fu_LIFTING_U3 ( .A(fu_LIFTING_n83), .Y(fu_LIFTING_n1) );
  DFFSX2 fu_LIFTING_reg_out_reg_31_ ( .D(fu_LIFTING_n442), .CK(clk), .SN(rstx), 
        .QN(ic_socket_LIFTING_o1_data0_wire[31]) );
  DFFSX2 fu_LIFTING_reg_out_reg_30_ ( .D(fu_LIFTING_n441), .CK(clk), .SN(rstx), 
        .QN(ic_socket_LIFTING_o1_data0_wire[30]) );
  DFFSX2 fu_LIFTING_reg_out_reg_29_ ( .D(fu_LIFTING_n440), .CK(clk), .SN(rstx), 
        .QN(ic_socket_LIFTING_o1_data0_wire[29]) );
  DFFSX2 fu_LIFTING_reg_out_reg_28_ ( .D(fu_LIFTING_n439), .CK(clk), .SN(rstx), 
        .QN(ic_socket_LIFTING_o1_data0_wire[28]) );
  DFFSX2 fu_LIFTING_reg_out_reg_27_ ( .D(fu_LIFTING_n438), .CK(clk), .SN(rstx), 
        .QN(ic_socket_LIFTING_o1_data0_wire[27]) );
  DFFSX2 fu_LIFTING_reg_out_reg_26_ ( .D(fu_LIFTING_n437), .CK(clk), .SN(rstx), 
        .QN(ic_socket_LIFTING_o1_data0_wire[26]) );
  DFFSX2 fu_LIFTING_reg_out_reg_25_ ( .D(fu_LIFTING_n436), .CK(clk), .SN(rstx), 
        .QN(ic_socket_LIFTING_o1_data0_wire[25]) );
  DFFSX2 fu_LIFTING_reg_out_reg_24_ ( .D(fu_LIFTING_n435), .CK(clk), .SN(rstx), 
        .QN(ic_socket_LIFTING_o1_data0_wire[24]) );
  DFFSX2 fu_LIFTING_reg_out_reg_23_ ( .D(fu_LIFTING_n434), .CK(clk), .SN(rstx), 
        .QN(ic_socket_LIFTING_o1_data0_wire[23]) );
  DFFSX2 fu_LIFTING_reg_out_reg_22_ ( .D(fu_LIFTING_n433), .CK(clk), .SN(rstx), 
        .QN(ic_socket_LIFTING_o1_data0_wire[22]) );
  DFFSX2 fu_LIFTING_reg_out_reg_21_ ( .D(fu_LIFTING_n432), .CK(clk), .SN(rstx), 
        .QN(ic_socket_LIFTING_o1_data0_wire[21]) );
  DFFSX2 fu_LIFTING_reg_out_reg_20_ ( .D(fu_LIFTING_n431), .CK(clk), .SN(rstx), 
        .QN(ic_socket_LIFTING_o1_data0_wire[20]) );
  DFFSX2 fu_LIFTING_reg_out_reg_19_ ( .D(fu_LIFTING_n430), .CK(clk), .SN(rstx), 
        .QN(ic_socket_LIFTING_o1_data0_wire[19]) );
  DFFSX2 fu_LIFTING_reg_out_reg_18_ ( .D(fu_LIFTING_n429), .CK(clk), .SN(rstx), 
        .QN(ic_socket_LIFTING_o1_data0_wire[18]) );
  DFFSX2 fu_LIFTING_reg_out_reg_17_ ( .D(fu_LIFTING_n428), .CK(clk), .SN(rstx), 
        .QN(ic_socket_LIFTING_o1_data0_wire[17]) );
  DFFSX2 fu_LIFTING_reg_out_reg_16_ ( .D(fu_LIFTING_n427), .CK(clk), .SN(rstx), 
        .QN(ic_socket_LIFTING_o1_data0_wire[16]) );
  DFFSX2 fu_LIFTING_reg_out_reg_15_ ( .D(fu_LIFTING_n426), .CK(clk), .SN(rstx), 
        .QN(ic_socket_LIFTING_o1_data0_wire[15]) );
  DFFSX2 fu_LIFTING_reg_out_reg_14_ ( .D(fu_LIFTING_n425), .CK(clk), .SN(rstx), 
        .QN(ic_socket_LIFTING_o1_data0_wire[14]) );
  DFFSX2 fu_LIFTING_reg_out_reg_13_ ( .D(fu_LIFTING_n424), .CK(clk), .SN(rstx), 
        .QN(ic_socket_LIFTING_o1_data0_wire[13]) );
  DFFSX2 fu_LIFTING_reg_out_reg_12_ ( .D(fu_LIFTING_n423), .CK(clk), .SN(rstx), 
        .QN(ic_socket_LIFTING_o1_data0_wire[12]) );
  DFFSX2 fu_LIFTING_reg_out_reg_11_ ( .D(fu_LIFTING_n422), .CK(clk), .SN(rstx), 
        .QN(ic_socket_LIFTING_o1_data0_wire[11]) );
  DFFSX2 fu_LIFTING_reg_out_reg_10_ ( .D(fu_LIFTING_n421), .CK(clk), .SN(rstx), 
        .QN(ic_socket_LIFTING_o1_data0_wire[10]) );
  DFFSX2 fu_LIFTING_reg_out_reg_9_ ( .D(fu_LIFTING_n420), .CK(clk), .SN(rstx), 
        .QN(ic_socket_LIFTING_o1_data0_wire[9]) );
  DFFSX2 fu_LIFTING_reg_out_reg_8_ ( .D(fu_LIFTING_n419), .CK(clk), .SN(rstx), 
        .QN(ic_socket_LIFTING_o1_data0_wire[8]) );
  DFFSX2 fu_LIFTING_reg_out_reg_7_ ( .D(fu_LIFTING_n418), .CK(clk), .SN(rstx), 
        .QN(ic_socket_LIFTING_o1_data0_wire[7]) );
  DFFSX2 fu_LIFTING_reg_out_reg_6_ ( .D(fu_LIFTING_n417), .CK(clk), .SN(rstx), 
        .QN(ic_socket_LIFTING_o1_data0_wire[6]) );
  DFFSX2 fu_LIFTING_reg_out_reg_5_ ( .D(fu_LIFTING_n416), .CK(clk), .SN(rstx), 
        .QN(ic_socket_LIFTING_o1_data0_wire[5]) );
  DFFSX2 fu_LIFTING_reg_out_reg_4_ ( .D(fu_LIFTING_n415), .CK(clk), .SN(rstx), 
        .QN(ic_socket_LIFTING_o1_data0_wire[4]) );
  DFFSX2 fu_LIFTING_reg_out_reg_3_ ( .D(fu_LIFTING_n414), .CK(clk), .SN(rstx), 
        .QN(ic_socket_LIFTING_o1_data0_wire[3]) );
  DFFSX2 fu_LIFTING_reg_out_reg_2_ ( .D(fu_LIFTING_n413), .CK(clk), .SN(rstx), 
        .QN(ic_socket_LIFTING_o1_data0_wire[2]) );
  DFFSX2 fu_LIFTING_reg_out_reg_1_ ( .D(fu_LIFTING_n412), .CK(clk), .SN(rstx), 
        .QN(ic_socket_LIFTING_o1_data0_wire[1]) );
  DFFSX2 fu_LIFTING_reg_out_reg_0_ ( .D(fu_LIFTING_n411), .CK(clk), .SN(rstx), 
        .QN(ic_socket_LIFTING_o1_data0_wire[0]) );
  CLKXOR2X2 fu_LIFTING_sub_98_DP_OP_282_1544_7_U50 ( .A(fu_LIFTING_n41), .B(
        fu_LIFTING_n496), .Y(fu_LIFTING_sub_98_DP_OP_282_1544_7_n51) );
  CLKXOR2X2 fu_LIFTING_sub_98_DP_OP_282_1544_7_U44 ( .A(fu_LIFTING_n41), .B(
        fu_LIFTING_n500), .Y(fu_LIFTING_sub_98_DP_OP_282_1544_7_n45) );
  CLKXOR2X2 fu_LIFTING_sub_98_DP_OP_282_1544_7_U41 ( .A(fu_LIFTING_n41), .B(
        fu_LIFTING_n500), .Y(fu_LIFTING_sub_98_DP_OP_282_1544_7_n42) );
  CLKXOR2X2 fu_LIFTING_sub_98_DP_OP_282_1544_7_U42 ( .A(fu_LIFTING_n41), .B(
        fu_LIFTING_n500), .Y(fu_LIFTING_sub_98_DP_OP_282_1544_7_n43) );
  CLKXOR2X2 fu_LIFTING_sub_98_DP_OP_282_1544_7_U43 ( .A(fu_LIFTING_n41), .B(
        fu_LIFTING_n500), .Y(fu_LIFTING_sub_98_DP_OP_282_1544_7_n44) );
  CLKXOR2X2 fu_LIFTING_sub_98_DP_OP_282_1544_7_U40 ( .A(fu_LIFTING_n41), .B(
        fu_LIFTING_n500), .Y(fu_LIFTING_sub_98_DP_OP_282_1544_7_n41) );
  CLKXOR2X2 fu_LIFTING_sub_98_DP_OP_282_1544_7_U39 ( .A(fu_LIFTING_n41), .B(
        fu_LIFTING_n500), .Y(fu_LIFTING_sub_98_DP_OP_282_1544_7_n40) );
  ADDFX2 fu_LIFTING_sub_98_DP_OP_282_1544_7_U17 ( .A(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n54), .B(fu_LIFTING_n459), .CI(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n17), .CO(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n16), .S(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_16_) );
  ADDFX2 fu_LIFTING_sub_98_DP_OP_282_1544_7_U18 ( .A(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n55), .B(fu_LIFTING_n458), .CI(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n18), .CO(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n17), .S(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_15_) );
  ADDFX2 fu_LIFTING_sub_98_DP_OP_282_1544_7_U19 ( .A(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n56), .B(fu_LIFTING_n457), .CI(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n19), .CO(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n18), .S(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_14_) );
  ADDFX1 fu_LIFTING_mult_84_DP_OP_276_6650_3_U32 ( .A(fu_LIFTING_N677), .B(
        fu_LIFTING_N673), .CI(fu_LIFTING_N676), .CO(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n31), .S(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n32) );
  ADDFX1 fu_LIFTING_mult_92_DP_OP_280_6650_5_U34 ( .A(fu_LIFTING_N679), .B(
        fu_LIFTING_n43), .CI(fu_LIFTING_N677), .CO(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n33), .S(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n34) );
  ADDFX1 fu_LIFTING_mult_84_DP_OP_276_6650_3_U33 ( .A(fu_LIFTING_N678), .B(
        fu_LIFTING_N674), .CI(fu_LIFTING_N677), .CO(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n33), .S(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n34) );
  ADDFX1 fu_LIFTING_mult_96_DP_OP_281_6650_6_U35 ( .A(fu_LIFTING_N81), .B(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n83), .CI(fu_LIFTING_N78), .CO(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n35), .S(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n36) );
  ADDFX1 fu_LIFTING_mult_92_DP_OP_280_6650_5_U35 ( .A(fu_LIFTING_N680), .B(
        fu_LIFTING_n44), .CI(fu_LIFTING_N678), .CO(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n35), .S(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n36) );
  ADDFX1 fu_LIFTING_mult_88_DP_OP_277_6650_4_U32 ( .A(fu_LIFTING_N79), .B(
        fu_LIFTING_N75), .CI(fu_LIFTING_N78), .CO(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n32), .S(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n33) );
  ADDFX4 fu_LIFTING_mult_96_DP_OP_281_6650_6_U4 ( .A(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n36), .B(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n37), .CI(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n4), .CO(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n3), .S(fu_LIFTING_N669) );
  ADDFX2 fu_LIFTING_sub_98_DP_OP_282_1544_7_U20 ( .A(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n57), .B(fu_LIFTING_n456), .CI(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n20), .CO(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n19), .S(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_13_) );
  ADDFX2 fu_LIFTING_sub_98_DP_OP_282_1544_7_U21 ( .A(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n58), .B(fu_LIFTING_n455), .CI(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n21), .CO(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n20), .S(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_12_) );
  ADDFX2 fu_LIFTING_sub_98_DP_OP_282_1544_7_U22 ( .A(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n59), .B(fu_LIFTING_n454), .CI(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n22), .CO(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n21), .S(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_11_) );
  ADDFX2 fu_LIFTING_mult_88_DP_OP_277_6650_4_U7 ( .A(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n39), .B(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n40), .CI(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n7), .CO(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n6), .S(fu_LIFTING_N426) );
  ADDFX2 fu_LIFTING_mult_79_DP_OP_279_6650_2_U6 ( .A(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n36), .B(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n37), .CI(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n6), .CO(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n5), .S(fu_LIFTING_N187) );
  ADDFX1 fu_LIFTING_mult_96_DP_OP_281_6650_6_U34 ( .A(fu_LIFTING_N80), .B(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n82), .CI(fu_LIFTING_N77), .CO(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n33), .S(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n34) );
  ADDFX1 fu_LIFTING_mult_88_DP_OP_277_6650_4_U31 ( .A(fu_LIFTING_N78), .B(
        fu_LIFTING_N74), .CI(fu_LIFTING_N77), .CO(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n30), .S(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n31) );
  ADDFX1 fu_LIFTING_mult_79_DP_OP_279_6650_2_U30 ( .A(fu_LIFTING_N79), .B(
        fu_LIFTING_N74), .CI(fu_LIFTING_N78), .CO(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n29), .S(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n30) );
  ADDFX1 fu_LIFTING_mult_79_DP_OP_279_6650_2_U31 ( .A(fu_LIFTING_N80), .B(
        fu_LIFTING_N75), .CI(fu_LIFTING_N79), .CO(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n31), .S(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n32) );
  CLKXOR2X2 fu_LIFTING_sub_98_DP_OP_282_1544_7_U2 ( .A(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n39), .B(fu_LIFTING_n474), .Y(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n1) );
  CLKXOR2X2 fu_LIFTING_sub_98_DP_OP_282_1544_7_U38 ( .A(fu_LIFTING_n41), .B(
        fu_LIFTING_n500), .Y(fu_LIFTING_sub_98_DP_OP_282_1544_7_n39) );
  ADDFX2 fu_LIFTING_mult_96_DP_OP_281_6650_6_U7 ( .A(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n42), .B(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n43), .CI(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n7), .CO(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n6), .S(fu_LIFTING_N666) );
  ADDFX2 fu_LIFTING_mult_96_DP_OP_281_6650_6_U8 ( .A(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n44), .B(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n45), .CI(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n8), .CO(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n7), .S(fu_LIFTING_N665) );
  ADDFX2 fu_LIFTING_mult_88_DP_OP_277_6650_4_U6 ( .A(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n37), .B(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n38), .CI(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n6), .CO(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n5), .S(fu_LIFTING_N427) );
  ADDFX2 fu_LIFTING_sub_98_DP_OP_282_1544_7_U23 ( .A(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n60), .B(fu_LIFTING_n453), .CI(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n23), .CO(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n22), .S(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_10_) );
  OR2X2 fu_LIFTING_sub_98_DP_OP_282_1544_7_U71 ( .A(fu_LIFTING_n238), .B(
        fu_LIFTING_n240), .Y(fu_LIFTING_sub_98_DP_OP_282_1544_7_n72) );
  NAND2X2 fu_LIFTING_U76 ( .A(fu_LIFTING_t1opcode_wire[2]), .B(
        fu_LIFTING_t1opcode_wire[1]), .Y(fu_LIFTING_n107) );
  CLKXOR2X2 fu_LIFTING_sub_98_DP_OP_282_1544_7_U59 ( .A(fu_LIFTING_n41), .B(
        fu_LIFTING_n487), .Y(fu_LIFTING_sub_98_DP_OP_282_1544_7_n60) );
  CLKXOR2X2 fu_LIFTING_sub_98_DP_OP_282_1544_7_U60 ( .A(fu_LIFTING_n41), .B(
        fu_LIFTING_n486), .Y(fu_LIFTING_sub_98_DP_OP_282_1544_7_n61) );
  CLKXOR2X2 fu_LIFTING_sub_98_DP_OP_282_1544_7_U61 ( .A(fu_LIFTING_n41), .B(
        fu_LIFTING_n485), .Y(fu_LIFTING_sub_98_DP_OP_282_1544_7_n62) );
  ADDFX4 fu_LIFTING_sub_98_DP_OP_282_1544_7_U4 ( .A(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n41), .B(fu_LIFTING_n472), .CI(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n4), .CO(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n3), .S(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_29_) );
  ADDFX4 fu_LIFTING_sub_98_DP_OP_282_1544_7_U12 ( .A(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n49), .B(fu_LIFTING_n464), .CI(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n12), .CO(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n11), .S(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_21_) );
  ADDFX4 fu_LIFTING_sub_98_DP_OP_282_1544_7_U13 ( .A(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n50), .B(fu_LIFTING_n463), .CI(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n13), .CO(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n12), .S(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_20_) );
  ADDFX4 fu_LIFTING_sub_98_DP_OP_282_1544_7_U16 ( .A(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n53), .B(fu_LIFTING_n460), .CI(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n16), .CO(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n15), .S(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_17_) );
  OR2X2 fu_LIFTING_sub_98_DP_OP_282_1544_7_U70 ( .A(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n72), .B(fu_LIFTING_n83), .Y(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n71) );
  CLKXOR2X2 fu_LIFTING_sub_98_DP_OP_282_1544_7_U56 ( .A(fu_LIFTING_n41), .B(
        fu_LIFTING_n490), .Y(fu_LIFTING_sub_98_DP_OP_282_1544_7_n57) );
  CLKXOR2X2 fu_LIFTING_sub_98_DP_OP_282_1544_7_U57 ( .A(fu_LIFTING_n41), .B(
        fu_LIFTING_n489), .Y(fu_LIFTING_sub_98_DP_OP_282_1544_7_n58) );
  CLKXOR2X2 fu_LIFTING_sub_98_DP_OP_282_1544_7_U58 ( .A(fu_LIFTING_n41), .B(
        fu_LIFTING_n488), .Y(fu_LIFTING_sub_98_DP_OP_282_1544_7_n59) );
  ADDFX2 fu_LIFTING_sub_98_DP_OP_282_1544_7_U24 ( .A(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n61), .B(fu_LIFTING_n452), .CI(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n24), .CO(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n23), .S(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_9_) );
  ADDFX4 fu_LIFTING_sub_98_DP_OP_282_1544_7_U5 ( .A(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n42), .B(fu_LIFTING_n471), .CI(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n5), .CO(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n4), .S(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_28_) );
  ADDFX4 fu_LIFTING_sub_98_DP_OP_282_1544_7_U6 ( .A(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n43), .B(fu_LIFTING_n470), .CI(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n6), .CO(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n5), .S(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_27_) );
  ADDFX4 fu_LIFTING_sub_98_DP_OP_282_1544_7_U7 ( .A(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n44), .B(fu_LIFTING_n469), .CI(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n7), .CO(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n6), .S(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_26_) );
  ADDFX2 fu_LIFTING_sub_98_DP_OP_282_1544_7_U25 ( .A(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n62), .B(fu_LIFTING_n451), .CI(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n25), .CO(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n24), .S(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_8_) );
  ADDFX2 fu_LIFTING_sub_98_DP_OP_282_1544_7_U26 ( .A(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n63), .B(fu_LIFTING_n450), .CI(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n26), .CO(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n25), .S(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_7_) );
  ADDFX2 fu_LIFTING_sub_98_DP_OP_282_1544_7_U27 ( .A(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n64), .B(fu_LIFTING_n449), .CI(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n27), .CO(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n26), .S(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_6_) );
  ADDFX2 fu_LIFTING_sub_98_DP_OP_282_1544_7_U28 ( .A(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n65), .B(fu_LIFTING_n448), .CI(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n28), .CO(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n27), .S(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_5_) );
  ADDFX2 fu_LIFTING_sub_98_DP_OP_282_1544_7_U29 ( .A(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n66), .B(fu_LIFTING_n447), .CI(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n29), .CO(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n28), .S(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_4_) );
  ADDFX2 fu_LIFTING_sub_98_DP_OP_282_1544_7_U30 ( .A(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n67), .B(fu_LIFTING_n446), .CI(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n30), .CO(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n29), .S(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_3_) );
  ADDFX2 fu_LIFTING_sub_98_DP_OP_282_1544_7_U31 ( .A(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n68), .B(fu_LIFTING_n445), .CI(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n31), .CO(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n30), .S(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_2_) );
  ADDFX2 fu_LIFTING_sub_98_DP_OP_282_1544_7_U32 ( .A(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n69), .B(fu_LIFTING_n444), .CI(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n32), .CO(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n31), .S(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_1_) );
  ADDFX2 fu_LIFTING_sub_98_DP_OP_282_1544_7_U33 ( .A(fu_LIFTING_n41), .B(
        fu_LIFTING_n443), .CI(fu_LIFTING_sub_98_DP_OP_282_1544_7_n70), .CO(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_n32), .S(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_0_) );
  CMPR42X1 fu_LIFTING_mult_75_DP_OP_278_6650_1_U37 ( .A(fu_LIFTING_N677), .B(
        fu_LIFTING_N678), .C(fu_LIFTING_N674), .D(fu_LIFTING_N673), .ICI(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n39), .S(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n38), .ICO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n36), .CO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n37) );
  CMPR42X1 fu_LIFTING_mult_75_DP_OP_278_6650_1_U38 ( .A(fu_LIFTING_N678), .B(
        fu_LIFTING_N679), .C(fu_LIFTING_N675), .D(fu_LIFTING_N674), .ICI(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n42), .S(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n41), .ICO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n39), .CO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n40) );
  CMPR42X1 fu_LIFTING_mult_75_DP_OP_278_6650_1_U39 ( .A(fu_LIFTING_N679), .B(
        fu_LIFTING_N680), .C(fu_LIFTING_N676), .D(fu_LIFTING_N675), .ICI(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n45), .S(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n44), .ICO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n42), .CO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n43) );
  CMPR42X1 fu_LIFTING_mult_75_DP_OP_278_6650_1_U40 ( .A(fu_LIFTING_N680), .B(
        fu_LIFTING_N681), .C(fu_LIFTING_N677), .D(fu_LIFTING_N676), .ICI(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n48), .S(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n47), .ICO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n45), .CO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n46) );
  CMPR42X1 fu_LIFTING_mult_75_DP_OP_278_6650_1_U41 ( .A(fu_LIFTING_N681), .B(
        fu_LIFTING_N682), .C(fu_LIFTING_N678), .D(fu_LIFTING_N677), .ICI(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n51), .S(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n50), .ICO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n48), .CO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n49) );
  CMPR42X1 fu_LIFTING_mult_75_DP_OP_278_6650_1_U42 ( .A(fu_LIFTING_N682), .B(
        fu_LIFTING_N683), .C(fu_LIFTING_N679), .D(fu_LIFTING_N678), .ICI(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n54), .S(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n53), .ICO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n51), .CO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n52) );
  CMPR42X1 fu_LIFTING_mult_75_DP_OP_278_6650_1_U43 ( .A(fu_LIFTING_N683), .B(
        fu_LIFTING_N684), .C(fu_LIFTING_N680), .D(fu_LIFTING_N679), .ICI(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n57), .S(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n56), .ICO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n54), .CO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n55) );
  CMPR42X1 fu_LIFTING_mult_75_DP_OP_278_6650_1_U44 ( .A(fu_LIFTING_N684), .B(
        fu_LIFTING_N685), .C(fu_LIFTING_N681), .D(fu_LIFTING_N680), .ICI(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n60), .S(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n59), .ICO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n57), .CO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n58) );
  CMPR42X1 fu_LIFTING_mult_75_DP_OP_278_6650_1_U45 ( .A(fu_LIFTING_N685), .B(
        fu_LIFTING_N686), .C(fu_LIFTING_N682), .D(fu_LIFTING_N681), .ICI(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n63), .S(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n62), .ICO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n60), .CO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n61) );
  CMPR42X1 fu_LIFTING_mult_75_DP_OP_278_6650_1_U46 ( .A(fu_LIFTING_N686), .B(
        fu_LIFTING_N687), .C(fu_LIFTING_N683), .D(fu_LIFTING_N682), .ICI(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n66), .S(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n65), .ICO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n63), .CO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n64) );
  CMPR42X1 fu_LIFTING_mult_75_DP_OP_278_6650_1_U49 ( .A(fu_LIFTING_N689), .B(
        fu_LIFTING_N690), .C(fu_LIFTING_N686), .D(fu_LIFTING_N685), .ICI(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n75), .S(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n74), .ICO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n72), .CO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n73) );
  CMPR42X1 fu_LIFTING_mult_75_DP_OP_278_6650_1_U50 ( .A(fu_LIFTING_N690), .B(
        fu_LIFTING_N691), .C(fu_LIFTING_N687), .D(fu_LIFTING_N686), .ICI(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n78), .S(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n77), .ICO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n75), .CO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n76) );
  CMPR42X1 fu_LIFTING_mult_75_DP_OP_278_6650_1_U51 ( .A(fu_LIFTING_N691), .B(
        fu_LIFTING_N692), .C(fu_LIFTING_N688), .D(fu_LIFTING_N687), .ICI(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n81), .S(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n80), .ICO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n78), .CO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n79) );
  CMPR42X1 fu_LIFTING_mult_75_DP_OP_278_6650_1_U52 ( .A(fu_LIFTING_N692), .B(
        fu_LIFTING_N693), .C(fu_LIFTING_N689), .D(fu_LIFTING_N688), .ICI(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n84), .S(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n83), .ICO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n81), .CO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n82) );
  CMPR42X1 fu_LIFTING_mult_75_DP_OP_278_6650_1_U53 ( .A(fu_LIFTING_N693), .B(
        fu_LIFTING_N694), .C(fu_LIFTING_N690), .D(fu_LIFTING_N689), .ICI(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n87), .S(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n86), .ICO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n84), .CO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n85) );
  CMPR42X1 fu_LIFTING_mult_75_DP_OP_278_6650_1_U54 ( .A(fu_LIFTING_N694), .B(
        fu_LIFTING_N695), .C(fu_LIFTING_N691), .D(fu_LIFTING_N690), .ICI(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n90), .S(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n89), .ICO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n87), .CO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n88) );
  CMPR42X1 fu_LIFTING_mult_75_DP_OP_278_6650_1_U55 ( .A(fu_LIFTING_N695), .B(
        fu_LIFTING_N696), .C(fu_LIFTING_N692), .D(fu_LIFTING_N691), .ICI(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n93), .S(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n92), .ICO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n90), .CO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n91) );
  CMPR42X1 fu_LIFTING_mult_75_DP_OP_278_6650_1_U56 ( .A(fu_LIFTING_N696), .B(
        fu_LIFTING_N697), .C(fu_LIFTING_N693), .D(fu_LIFTING_N692), .ICI(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n96), .S(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n95), .ICO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n93), .CO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n94) );
  CMPR42X1 fu_LIFTING_mult_75_DP_OP_278_6650_1_U57 ( .A(fu_LIFTING_N697), .B(
        fu_LIFTING_N698), .C(fu_LIFTING_N694), .D(fu_LIFTING_N693), .ICI(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n99), .S(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n98), .ICO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n96), .CO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n97) );
  CMPR42X1 fu_LIFTING_mult_75_DP_OP_278_6650_1_U58 ( .A(fu_LIFTING_N698), .B(
        fu_LIFTING_N699), .C(fu_LIFTING_N695), .D(fu_LIFTING_N694), .ICI(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n102), .S(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n101), .ICO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n99), .CO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n100) );
  CMPR42X1 fu_LIFTING_mult_75_DP_OP_278_6650_1_U59 ( .A(fu_LIFTING_N699), .B(
        fu_LIFTING_N700), .C(fu_LIFTING_N696), .D(fu_LIFTING_N695), .ICI(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n105), .S(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n104), .ICO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n102), .CO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n103) );
  CMPR42X1 fu_LIFTING_mult_75_DP_OP_278_6650_1_U60 ( .A(fu_LIFTING_N700), .B(
        fu_LIFTING_N701), .C(fu_LIFTING_N697), .D(fu_LIFTING_N696), .ICI(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n108), .S(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n107), .ICO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n105), .CO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n106) );
  CMPR42X1 fu_LIFTING_mult_75_DP_OP_278_6650_1_U61 ( .A(fu_LIFTING_N701), .B(
        fu_LIFTING_N702), .C(fu_LIFTING_N698), .D(fu_LIFTING_N697), .ICI(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n113), .S(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n110), .ICO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n108), .CO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n109) );
  ADDFX2 fu_LIFTING_mult_75_DP_OP_278_6650_1_U4 ( .A(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n41), .B(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n43), .CI(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n4), .CO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n3), .S(fu_LIFTING_N69) );
  ADDFX2 fu_LIFTING_mult_75_DP_OP_278_6650_1_U7 ( .A(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n50), .B(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n52), .CI(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n7), .CO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n6), .S(fu_LIFTING_N66) );
  ADDFX1 fu_LIFTING_mult_75_DP_OP_278_6650_1_U8 ( .A(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n53), .B(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n55), .CI(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n8), .CO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n7), .S(fu_LIFTING_N65) );
  ADDFX1 fu_LIFTING_mult_75_DP_OP_278_6650_1_U16 ( .A(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n77), .B(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n79), .CI(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n16), .CO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n15), .S(fu_LIFTING_N57) );
  ADDFX1 fu_LIFTING_mult_75_DP_OP_278_6650_1_U17 ( .A(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n80), .B(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n82), .CI(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n17), .CO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n16), .S(fu_LIFTING_N56) );
  ADDFX1 fu_LIFTING_mult_75_DP_OP_278_6650_1_U18 ( .A(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n83), .B(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n85), .CI(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n18), .CO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n17), .S(fu_LIFTING_N55) );
  ADDFX1 fu_LIFTING_mult_75_DP_OP_278_6650_1_U19 ( .A(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n86), .B(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n88), .CI(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n19), .CO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n18), .S(fu_LIFTING_N54) );
  ADDFX1 fu_LIFTING_mult_75_DP_OP_278_6650_1_U25 ( .A(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n104), .B(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n106), .CI(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n25), .CO(
        fu_LIFTING_mult_75_DP_OP_278_6650_1_n24), .S(fu_LIFTING_N48) );
  ADDFX1 fu_LIFTING_mult_79_DP_OP_279_6650_2_U33 ( .A(fu_LIFTING_N82), .B(
        fu_LIFTING_N77), .CI(fu_LIFTING_N81), .CO(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n35), .S(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n36) );
  ADDFX1 fu_LIFTING_mult_79_DP_OP_279_6650_2_U34 ( .A(fu_LIFTING_N83), .B(
        fu_LIFTING_N78), .CI(fu_LIFTING_N82), .CO(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n37), .S(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n38) );
  ADDFX1 fu_LIFTING_mult_79_DP_OP_279_6650_2_U35 ( .A(fu_LIFTING_N84), .B(
        fu_LIFTING_N79), .CI(fu_LIFTING_N83), .CO(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n39), .S(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n40) );
  ADDFX1 fu_LIFTING_mult_79_DP_OP_279_6650_2_U36 ( .A(fu_LIFTING_N85), .B(
        fu_LIFTING_N80), .CI(fu_LIFTING_N84), .CO(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n41), .S(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n42) );
  ADDFX1 fu_LIFTING_mult_79_DP_OP_279_6650_2_U37 ( .A(fu_LIFTING_N86), .B(
        fu_LIFTING_N81), .CI(fu_LIFTING_N85), .CO(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n43), .S(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n44) );
  ADDFX1 fu_LIFTING_mult_79_DP_OP_279_6650_2_U38 ( .A(fu_LIFTING_N87), .B(
        fu_LIFTING_N82), .CI(fu_LIFTING_N86), .CO(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n45), .S(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n46) );
  ADDFX1 fu_LIFTING_mult_79_DP_OP_279_6650_2_U39 ( .A(fu_LIFTING_N88), .B(
        fu_LIFTING_N83), .CI(fu_LIFTING_N87), .CO(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n47), .S(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n48) );
  ADDFX1 fu_LIFTING_mult_79_DP_OP_279_6650_2_U40 ( .A(fu_LIFTING_N89), .B(
        fu_LIFTING_N84), .CI(fu_LIFTING_N88), .CO(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n49), .S(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n50) );
  ADDFX1 fu_LIFTING_mult_79_DP_OP_279_6650_2_U42 ( .A(fu_LIFTING_N91), .B(
        fu_LIFTING_N86), .CI(fu_LIFTING_N90), .CO(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n53), .S(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n54) );
  ADDFX1 fu_LIFTING_mult_79_DP_OP_279_6650_2_U44 ( .A(fu_LIFTING_N93), .B(
        fu_LIFTING_N88), .CI(fu_LIFTING_N92), .CO(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n57), .S(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n58) );
  ADDFX1 fu_LIFTING_mult_79_DP_OP_279_6650_2_U45 ( .A(fu_LIFTING_N94), .B(
        fu_LIFTING_N89), .CI(fu_LIFTING_N93), .CO(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n59), .S(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n60) );
  ADDFX1 fu_LIFTING_mult_79_DP_OP_279_6650_2_U48 ( .A(fu_LIFTING_N97), .B(
        fu_LIFTING_N92), .CI(fu_LIFTING_N96), .CO(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n65), .S(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n66) );
  ADDFX1 fu_LIFTING_mult_79_DP_OP_279_6650_2_U49 ( .A(fu_LIFTING_N98), .B(
        fu_LIFTING_N93), .CI(fu_LIFTING_N97), .CO(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n67), .S(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n68) );
  ADDFX1 fu_LIFTING_mult_79_DP_OP_279_6650_2_U50 ( .A(fu_LIFTING_N99), .B(
        fu_LIFTING_N94), .CI(fu_LIFTING_N98), .CO(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n69), .S(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n70) );
  ADDFX1 fu_LIFTING_mult_79_DP_OP_279_6650_2_U25 ( .A(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n74), .B(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n75), .CI(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n25), .CO(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n24), .S(fu_LIFTING_N168) );
  ADDFX1 fu_LIFTING_mult_79_DP_OP_279_6650_2_U24 ( .A(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n72), .B(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n73), .CI(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n24), .CO(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n23), .S(fu_LIFTING_N169) );
  ADDFX1 fu_LIFTING_mult_79_DP_OP_279_6650_2_U23 ( .A(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n70), .B(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n71), .CI(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n23), .CO(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n22), .S(fu_LIFTING_N170) );
  ADDFX1 fu_LIFTING_mult_79_DP_OP_279_6650_2_U22 ( .A(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n68), .B(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n69), .CI(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n22), .CO(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n21), .S(fu_LIFTING_N171) );
  ADDFX1 fu_LIFTING_mult_79_DP_OP_279_6650_2_U21 ( .A(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n66), .B(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n67), .CI(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n21), .CO(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n20), .S(fu_LIFTING_N172) );
  ADDFX1 fu_LIFTING_mult_79_DP_OP_279_6650_2_U17 ( .A(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n58), .B(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n59), .CI(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n17), .CO(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n16), .S(fu_LIFTING_N176) );
  ADDFX1 fu_LIFTING_mult_79_DP_OP_279_6650_2_U7 ( .A(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n38), .B(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n39), .CI(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n7), .CO(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n6), .S(fu_LIFTING_N186) );
  ADDFX1 fu_LIFTING_mult_79_DP_OP_279_6650_2_U8 ( .A(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n40), .B(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n41), .CI(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n8), .CO(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n7), .S(fu_LIFTING_N185) );
  ADDFX1 fu_LIFTING_mult_79_DP_OP_279_6650_2_U11 ( .A(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n46), .B(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n47), .CI(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n11), .CO(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n10), .S(fu_LIFTING_N182) );
  ADDFX1 fu_LIFTING_mult_79_DP_OP_279_6650_2_U12 ( .A(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n48), .B(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n49), .CI(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n12), .CO(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n11), .S(fu_LIFTING_N181) );
  ADDFX1 fu_LIFTING_mult_79_DP_OP_279_6650_2_U16 ( .A(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n56), .B(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n57), .CI(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n16), .CO(
        fu_LIFTING_mult_79_DP_OP_279_6650_2_n15), .S(fu_LIFTING_N177) );
  ADDFX1 fu_LIFTING_mult_84_DP_OP_276_6650_3_U35 ( .A(fu_LIFTING_N680), .B(
        fu_LIFTING_N676), .CI(fu_LIFTING_N679), .CO(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n37), .S(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n38) );
  ADDFX1 fu_LIFTING_mult_84_DP_OP_276_6650_3_U37 ( .A(fu_LIFTING_N682), .B(
        fu_LIFTING_N678), .CI(fu_LIFTING_N681), .CO(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n41), .S(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n42) );
  ADDFX1 fu_LIFTING_mult_84_DP_OP_276_6650_3_U38 ( .A(fu_LIFTING_N683), .B(
        fu_LIFTING_N679), .CI(fu_LIFTING_N682), .CO(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n43), .S(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n44) );
  ADDFX1 fu_LIFTING_mult_84_DP_OP_276_6650_3_U39 ( .A(fu_LIFTING_N684), .B(
        fu_LIFTING_N680), .CI(fu_LIFTING_N683), .CO(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n45), .S(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n46) );
  ADDFX1 fu_LIFTING_mult_84_DP_OP_276_6650_3_U40 ( .A(fu_LIFTING_N685), .B(
        fu_LIFTING_N681), .CI(fu_LIFTING_N684), .CO(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n47), .S(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n48) );
  ADDFX1 fu_LIFTING_mult_84_DP_OP_276_6650_3_U41 ( .A(fu_LIFTING_N686), .B(
        fu_LIFTING_N682), .CI(fu_LIFTING_N685), .CO(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n49), .S(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n50) );
  ADDFX1 fu_LIFTING_mult_84_DP_OP_276_6650_3_U43 ( .A(fu_LIFTING_N688), .B(
        fu_LIFTING_N684), .CI(fu_LIFTING_N687), .CO(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n53), .S(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n54) );
  ADDFX1 fu_LIFTING_mult_84_DP_OP_276_6650_3_U44 ( .A(fu_LIFTING_N689), .B(
        fu_LIFTING_N685), .CI(fu_LIFTING_N688), .CO(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n55), .S(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n56) );
  ADDFX1 fu_LIFTING_mult_84_DP_OP_276_6650_3_U45 ( .A(fu_LIFTING_N690), .B(
        fu_LIFTING_N686), .CI(fu_LIFTING_N689), .CO(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n57), .S(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n58) );
  ADDFX1 fu_LIFTING_mult_84_DP_OP_276_6650_3_U46 ( .A(fu_LIFTING_N691), .B(
        fu_LIFTING_N687), .CI(fu_LIFTING_N690), .CO(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n59), .S(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n60) );
  ADDFX1 fu_LIFTING_mult_84_DP_OP_276_6650_3_U47 ( .A(fu_LIFTING_N692), .B(
        fu_LIFTING_N688), .CI(fu_LIFTING_N691), .CO(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n61), .S(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n62) );
  ADDFX1 fu_LIFTING_mult_84_DP_OP_276_6650_3_U48 ( .A(fu_LIFTING_N693), .B(
        fu_LIFTING_N689), .CI(fu_LIFTING_N692), .CO(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n63), .S(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n64) );
  ADDFX1 fu_LIFTING_mult_84_DP_OP_276_6650_3_U49 ( .A(fu_LIFTING_N694), .B(
        fu_LIFTING_N690), .CI(fu_LIFTING_N693), .CO(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n65), .S(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n66) );
  ADDFX1 fu_LIFTING_mult_84_DP_OP_276_6650_3_U50 ( .A(fu_LIFTING_N695), .B(
        fu_LIFTING_N691), .CI(fu_LIFTING_N694), .CO(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n67), .S(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n68) );
  ADDFX1 fu_LIFTING_mult_84_DP_OP_276_6650_3_U51 ( .A(fu_LIFTING_N696), .B(
        fu_LIFTING_N692), .CI(fu_LIFTING_N695), .CO(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n69), .S(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n70) );
  ADDFX1 fu_LIFTING_mult_84_DP_OP_276_6650_3_U52 ( .A(fu_LIFTING_N697), .B(
        fu_LIFTING_N693), .CI(fu_LIFTING_N696), .CO(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n71), .S(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n72) );
  ADDFX1 fu_LIFTING_mult_84_DP_OP_276_6650_3_U53 ( .A(fu_LIFTING_N698), .B(
        fu_LIFTING_N694), .CI(fu_LIFTING_N697), .CO(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n73), .S(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n74) );
  ADDFX1 fu_LIFTING_mult_84_DP_OP_276_6650_3_U54 ( .A(fu_LIFTING_N699), .B(
        fu_LIFTING_N695), .CI(fu_LIFTING_N698), .CO(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n75), .S(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n76) );
  ADDFX1 fu_LIFTING_mult_84_DP_OP_276_6650_3_U55 ( .A(fu_LIFTING_N700), .B(
        fu_LIFTING_N696), .CI(fu_LIFTING_N699), .CO(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n77), .S(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n78) );
  ADDFX1 fu_LIFTING_mult_84_DP_OP_276_6650_3_U34 ( .A(fu_LIFTING_N679), .B(
        fu_LIFTING_N675), .CI(fu_LIFTING_N678), .CO(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n35), .S(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n36) );
  ADDFX1 fu_LIFTING_mult_84_DP_OP_276_6650_3_U9 ( .A(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n44), .B(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n45), .CI(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n9), .CO(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n8), .S(fu_LIFTING_N304) );
  ADDFX1 fu_LIFTING_mult_84_DP_OP_276_6650_3_U10 ( .A(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n46), .B(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n47), .CI(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n10), .CO(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n9), .S(fu_LIFTING_N303) );
  ADDFX1 fu_LIFTING_mult_84_DP_OP_276_6650_3_U11 ( .A(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n48), .B(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n49), .CI(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n11), .CO(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n10), .S(fu_LIFTING_N302) );
  ADDFX1 fu_LIFTING_mult_84_DP_OP_276_6650_3_U18 ( .A(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n62), .B(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n63), .CI(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n18), .CO(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n17), .S(fu_LIFTING_N295) );
  ADDFX1 fu_LIFTING_mult_84_DP_OP_276_6650_3_U19 ( .A(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n64), .B(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n65), .CI(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n19), .CO(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n18), .S(fu_LIFTING_N294) );
  ADDFX1 fu_LIFTING_mult_84_DP_OP_276_6650_3_U20 ( .A(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n66), .B(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n67), .CI(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n20), .CO(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n19), .S(fu_LIFTING_N293) );
  ADDFX1 fu_LIFTING_mult_84_DP_OP_276_6650_3_U21 ( .A(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n68), .B(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n69), .CI(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n21), .CO(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n20), .S(fu_LIFTING_N292) );
  ADDFX1 fu_LIFTING_mult_84_DP_OP_276_6650_3_U25 ( .A(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n76), .B(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n77), .CI(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n25), .CO(
        fu_LIFTING_mult_84_DP_OP_276_6650_3_n24), .S(fu_LIFTING_N288) );
  ADDFX1 fu_LIFTING_mult_88_DP_OP_277_6650_4_U35 ( .A(fu_LIFTING_N82), .B(
        fu_LIFTING_N78), .CI(fu_LIFTING_N81), .CO(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n38), .S(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n39) );
  ADDFX1 fu_LIFTING_mult_88_DP_OP_277_6650_4_U36 ( .A(fu_LIFTING_N83), .B(
        fu_LIFTING_N79), .CI(fu_LIFTING_N82), .CO(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n40), .S(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n41) );
  ADDFX1 fu_LIFTING_mult_88_DP_OP_277_6650_4_U37 ( .A(fu_LIFTING_N84), .B(
        fu_LIFTING_N80), .CI(fu_LIFTING_N83), .CO(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n42), .S(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n43) );
  ADDFX1 fu_LIFTING_mult_88_DP_OP_277_6650_4_U38 ( .A(fu_LIFTING_N85), .B(
        fu_LIFTING_N81), .CI(fu_LIFTING_N84), .CO(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n44), .S(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n45) );
  ADDFX1 fu_LIFTING_mult_88_DP_OP_277_6650_4_U39 ( .A(fu_LIFTING_N86), .B(
        fu_LIFTING_N82), .CI(fu_LIFTING_N85), .CO(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n46), .S(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n47) );
  ADDFX1 fu_LIFTING_mult_88_DP_OP_277_6650_4_U40 ( .A(fu_LIFTING_N87), .B(
        fu_LIFTING_N83), .CI(fu_LIFTING_N86), .CO(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n48), .S(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n49) );
  ADDFX1 fu_LIFTING_mult_88_DP_OP_277_6650_4_U41 ( .A(fu_LIFTING_N88), .B(
        fu_LIFTING_N84), .CI(fu_LIFTING_N87), .CO(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n50), .S(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n51) );
  ADDFX1 fu_LIFTING_mult_88_DP_OP_277_6650_4_U43 ( .A(fu_LIFTING_N90), .B(
        fu_LIFTING_N86), .CI(fu_LIFTING_N89), .CO(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n54), .S(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n55) );
  ADDFX1 fu_LIFTING_mult_88_DP_OP_277_6650_4_U44 ( .A(fu_LIFTING_N91), .B(
        fu_LIFTING_N87), .CI(fu_LIFTING_N90), .CO(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n56), .S(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n57) );
  ADDFX1 fu_LIFTING_mult_88_DP_OP_277_6650_4_U45 ( .A(fu_LIFTING_N92), .B(
        fu_LIFTING_N88), .CI(fu_LIFTING_N91), .CO(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n58), .S(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n59) );
  ADDFX1 fu_LIFTING_mult_88_DP_OP_277_6650_4_U46 ( .A(fu_LIFTING_N93), .B(
        fu_LIFTING_N89), .CI(fu_LIFTING_N92), .CO(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n60), .S(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n61) );
  ADDFX1 fu_LIFTING_mult_88_DP_OP_277_6650_4_U47 ( .A(fu_LIFTING_N94), .B(
        fu_LIFTING_N90), .CI(fu_LIFTING_N93), .CO(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n62), .S(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n63) );
  ADDFX1 fu_LIFTING_mult_88_DP_OP_277_6650_4_U48 ( .A(fu_LIFTING_N95), .B(
        fu_LIFTING_N91), .CI(fu_LIFTING_N94), .CO(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n64), .S(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n65) );
  ADDFX1 fu_LIFTING_mult_88_DP_OP_277_6650_4_U8 ( .A(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n41), .B(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n42), .CI(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n8), .CO(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n7), .S(fu_LIFTING_N425) );
  ADDFX1 fu_LIFTING_mult_88_DP_OP_277_6650_4_U10 ( .A(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n45), .B(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n46), .CI(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n10), .CO(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n9), .S(fu_LIFTING_N423) );
  ADDFX1 fu_LIFTING_mult_88_DP_OP_277_6650_4_U11 ( .A(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n47), .B(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n48), .CI(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n11), .CO(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n10), .S(fu_LIFTING_N422) );
  ADDFX1 fu_LIFTING_mult_88_DP_OP_277_6650_4_U15 ( .A(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n55), .B(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n56), .CI(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n15), .CO(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n14), .S(fu_LIFTING_N418) );
  ADDFX1 fu_LIFTING_mult_88_DP_OP_277_6650_4_U16 ( .A(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n57), .B(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n58), .CI(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n16), .CO(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n15), .S(fu_LIFTING_N417) );
  ADDFX1 fu_LIFTING_mult_88_DP_OP_277_6650_4_U17 ( .A(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n59), .B(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n60), .CI(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n17), .CO(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n16), .S(fu_LIFTING_N416) );
  ADDFX1 fu_LIFTING_mult_88_DP_OP_277_6650_4_U18 ( .A(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n61), .B(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n62), .CI(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n18), .CO(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n17), .S(fu_LIFTING_N415) );
  ADDFX1 fu_LIFTING_mult_88_DP_OP_277_6650_4_U19 ( .A(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n63), .B(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n64), .CI(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n19), .CO(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n18), .S(fu_LIFTING_N414) );
  ADDFX1 fu_LIFTING_mult_88_DP_OP_277_6650_4_U20 ( .A(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n65), .B(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n66), .CI(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n20), .CO(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n19), .S(fu_LIFTING_N413) );
  ADDFX1 fu_LIFTING_mult_88_DP_OP_277_6650_4_U24 ( .A(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n73), .B(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n74), .CI(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n24), .CO(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n23), .S(fu_LIFTING_N409) );
  ADDFX1 fu_LIFTING_mult_88_DP_OP_277_6650_4_U25 ( .A(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n75), .B(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n76), .CI(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n25), .CO(
        fu_LIFTING_mult_88_DP_OP_277_6650_4_n24), .S(fu_LIFTING_N408) );
  ADDFX1 fu_LIFTING_mult_92_DP_OP_280_6650_5_U36 ( .A(fu_LIFTING_N681), .B(
        fu_LIFTING_n46), .CI(fu_LIFTING_N679), .CO(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n37), .S(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n38) );
  ADDFX1 fu_LIFTING_mult_92_DP_OP_280_6650_5_U37 ( .A(fu_LIFTING_N682), .B(
        fu_LIFTING_n47), .CI(fu_LIFTING_N680), .CO(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n39), .S(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n40) );
  ADDFX1 fu_LIFTING_mult_92_DP_OP_280_6650_5_U38 ( .A(fu_LIFTING_N683), .B(
        fu_LIFTING_n49), .CI(fu_LIFTING_N681), .CO(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n41), .S(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n42) );
  ADDFX1 fu_LIFTING_mult_92_DP_OP_280_6650_5_U39 ( .A(fu_LIFTING_N684), .B(
        fu_LIFTING_n50), .CI(fu_LIFTING_N682), .CO(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n43), .S(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n44) );
  ADDFX1 fu_LIFTING_mult_92_DP_OP_280_6650_5_U40 ( .A(fu_LIFTING_N685), .B(
        fu_LIFTING_n52), .CI(fu_LIFTING_N683), .CO(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n45), .S(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n46) );
  ADDFX1 fu_LIFTING_mult_92_DP_OP_280_6650_5_U41 ( .A(fu_LIFTING_N686), .B(
        fu_LIFTING_n53), .CI(fu_LIFTING_N684), .CO(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n47), .S(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n48) );
  ADDFX1 fu_LIFTING_mult_92_DP_OP_280_6650_5_U42 ( .A(fu_LIFTING_N687), .B(
        fu_LIFTING_n54), .CI(fu_LIFTING_N685), .CO(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n49), .S(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n50) );
  ADDFX1 fu_LIFTING_mult_92_DP_OP_280_6650_5_U43 ( .A(fu_LIFTING_N688), .B(
        fu_LIFTING_n55), .CI(fu_LIFTING_N686), .CO(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n51), .S(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n52) );
  ADDFX1 fu_LIFTING_mult_92_DP_OP_280_6650_5_U46 ( .A(fu_LIFTING_N691), .B(
        fu_LIFTING_n59), .CI(fu_LIFTING_N689), .CO(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n57), .S(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n58) );
  ADDFX1 fu_LIFTING_mult_92_DP_OP_280_6650_5_U47 ( .A(fu_LIFTING_N692), .B(
        fu_LIFTING_n60), .CI(fu_LIFTING_N690), .CO(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n59), .S(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n60) );
  ADDFX1 fu_LIFTING_mult_92_DP_OP_280_6650_5_U48 ( .A(fu_LIFTING_N693), .B(
        fu_LIFTING_n63), .CI(fu_LIFTING_N691), .CO(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n61), .S(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n62) );
  ADDFX1 fu_LIFTING_mult_92_DP_OP_280_6650_5_U49 ( .A(fu_LIFTING_N694), .B(
        fu_LIFTING_n61), .CI(fu_LIFTING_N692), .CO(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n63), .S(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n64) );
  ADDFX1 fu_LIFTING_mult_92_DP_OP_280_6650_5_U50 ( .A(fu_LIFTING_N695), .B(
        fu_LIFTING_n64), .CI(fu_LIFTING_N693), .CO(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n65), .S(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n66) );
  ADDFX1 fu_LIFTING_mult_92_DP_OP_280_6650_5_U51 ( .A(fu_LIFTING_N696), .B(
        fu_LIFTING_n66), .CI(fu_LIFTING_N694), .CO(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n67), .S(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n68) );
  ADDFX1 fu_LIFTING_mult_92_DP_OP_280_6650_5_U52 ( .A(fu_LIFTING_N697), .B(
        fu_LIFTING_n67), .CI(fu_LIFTING_N695), .CO(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n69), .S(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n70) );
  ADDFX1 fu_LIFTING_mult_92_DP_OP_280_6650_5_U55 ( .A(fu_LIFTING_N700), .B(
        fu_LIFTING_n81), .CI(fu_LIFTING_N698), .CO(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n75), .S(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n76) );
  ADDFX1 fu_LIFTING_mult_92_DP_OP_280_6650_5_U56 ( .A(fu_LIFTING_N701), .B(
        fu_LIFTING_n82), .CI(fu_LIFTING_N699), .CO(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n77), .S(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n78) );
  ADDFX1 fu_LIFTING_mult_92_DP_OP_280_6650_5_U57 ( .A(fu_LIFTING_N702), .B(
        fu_LIFTING_n80), .CI(fu_LIFTING_N700), .CO(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n79), .S(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n80) );
  ADDFX1 fu_LIFTING_mult_92_DP_OP_280_6650_5_U7 ( .A(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n42), .B(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n43), .CI(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n7), .CO(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n6), .S(fu_LIFTING_N546) );
  ADDFX1 fu_LIFTING_mult_92_DP_OP_280_6650_5_U15 ( .A(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n58), .B(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n59), .CI(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n15), .CO(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n14), .S(fu_LIFTING_N538) );
  ADDFX1 fu_LIFTING_mult_92_DP_OP_280_6650_5_U16 ( .A(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n60), .B(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n61), .CI(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n16), .CO(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n15), .S(fu_LIFTING_N537) );
  ADDFX1 fu_LIFTING_mult_92_DP_OP_280_6650_5_U17 ( .A(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n62), .B(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n63), .CI(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n17), .CO(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n16), .S(fu_LIFTING_N536) );
  ADDFX1 fu_LIFTING_mult_92_DP_OP_280_6650_5_U18 ( .A(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n64), .B(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n65), .CI(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n18), .CO(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n17), .S(fu_LIFTING_N535) );
  ADDFX1 fu_LIFTING_mult_92_DP_OP_280_6650_5_U20 ( .A(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n68), .B(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n69), .CI(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n20), .CO(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n19), .S(fu_LIFTING_N533) );
  ADDFX1 fu_LIFTING_mult_92_DP_OP_280_6650_5_U24 ( .A(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n76), .B(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n77), .CI(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n24), .CO(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n23), .S(fu_LIFTING_N529) );
  ADDFX1 fu_LIFTING_mult_92_DP_OP_280_6650_5_U25 ( .A(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n78), .B(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n79), .CI(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n25), .CO(
        fu_LIFTING_mult_92_DP_OP_280_6650_5_n24), .S(fu_LIFTING_N528) );
  ADDFX1 fu_LIFTING_mult_96_DP_OP_281_6650_6_U36 ( .A(fu_LIFTING_N82), .B(
        fu_LIFTING_n45), .CI(fu_LIFTING_N79), .CO(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n37), .S(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n38) );
  ADDFX1 fu_LIFTING_mult_96_DP_OP_281_6650_6_U39 ( .A(fu_LIFTING_N85), .B(
        fu_LIFTING_n51), .CI(fu_LIFTING_N82), .CO(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n43), .S(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n44) );
  ADDFX1 fu_LIFTING_mult_96_DP_OP_281_6650_6_U40 ( .A(fu_LIFTING_N86), .B(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n88), .CI(fu_LIFTING_N83), .CO(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n45), .S(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n46) );
  ADDFX1 fu_LIFTING_mult_96_DP_OP_281_6650_6_U41 ( .A(fu_LIFTING_N87), .B(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n89), .CI(fu_LIFTING_N84), .CO(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n47), .S(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n48) );
  ADDFX1 fu_LIFTING_mult_96_DP_OP_281_6650_6_U42 ( .A(fu_LIFTING_N88), .B(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n90), .CI(fu_LIFTING_N85), .CO(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n49), .S(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n50) );
  ADDFX1 fu_LIFTING_mult_96_DP_OP_281_6650_6_U43 ( .A(fu_LIFTING_N89), .B(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n91), .CI(fu_LIFTING_N86), .CO(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n51), .S(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n52) );
  ADDFX1 fu_LIFTING_mult_96_DP_OP_281_6650_6_U44 ( .A(fu_LIFTING_N90), .B(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n92), .CI(fu_LIFTING_N87), .CO(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n53), .S(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n54) );
  ADDFX1 fu_LIFTING_mult_96_DP_OP_281_6650_6_U45 ( .A(fu_LIFTING_N91), .B(
        fu_LIFTING_n58), .CI(fu_LIFTING_N88), .CO(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n55), .S(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n56) );
  ADDFX1 fu_LIFTING_mult_96_DP_OP_281_6650_6_U46 ( .A(fu_LIFTING_N92), .B(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n94), .CI(fu_LIFTING_N89), .CO(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n57), .S(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n58) );
  ADDFX1 fu_LIFTING_mult_96_DP_OP_281_6650_6_U49 ( .A(fu_LIFTING_N95), .B(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n97), .CI(fu_LIFTING_N92), .CO(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n63), .S(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n64) );
  ADDFX1 fu_LIFTING_mult_96_DP_OP_281_6650_6_U50 ( .A(fu_LIFTING_N96), .B(
        fu_LIFTING_n65), .CI(fu_LIFTING_N93), .CO(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n65), .S(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n66) );
  ADDFX1 fu_LIFTING_mult_96_DP_OP_281_6650_6_U51 ( .A(fu_LIFTING_N97), .B(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n99), .CI(fu_LIFTING_N94), .CO(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n67), .S(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n68) );
  ADDFX1 fu_LIFTING_mult_96_DP_OP_281_6650_6_U54 ( .A(fu_LIFTING_N644), .B(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n102), .CI(fu_LIFTING_N97), .CO(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n73), .S(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n74) );
  ADDFX1 fu_LIFTING_mult_96_DP_OP_281_6650_6_U55 ( .A(fu_LIFTING_N645), .B(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n103), .CI(fu_LIFTING_N98), .CO(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n75), .S(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n76) );
  ADDFX1 fu_LIFTING_mult_96_DP_OP_281_6650_6_U56 ( .A(fu_LIFTING_N646), .B(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n104), .CI(fu_LIFTING_N99), .CO(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n77), .S(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n78) );
  ADDFX1 fu_LIFTING_mult_96_DP_OP_281_6650_6_U9 ( .A(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n46), .B(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n47), .CI(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n9), .CO(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n8), .S(fu_LIFTING_N664) );
  ADDFX1 fu_LIFTING_mult_96_DP_OP_281_6650_6_U10 ( .A(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n48), .B(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n49), .CI(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n10), .CO(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n9), .S(fu_LIFTING_N663) );
  ADDFX1 fu_LIFTING_mult_96_DP_OP_281_6650_6_U14 ( .A(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n56), .B(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n57), .CI(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n14), .CO(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n13), .S(fu_LIFTING_N659) );
  ADDFX1 fu_LIFTING_mult_96_DP_OP_281_6650_6_U17 ( .A(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n62), .B(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n63), .CI(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n17), .CO(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n16), .S(fu_LIFTING_N656) );
  ADDFX1 fu_LIFTING_mult_96_DP_OP_281_6650_6_U18 ( .A(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n64), .B(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n65), .CI(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n18), .CO(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n17), .S(fu_LIFTING_N655) );
  ADDFX1 fu_LIFTING_mult_96_DP_OP_281_6650_6_U19 ( .A(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n66), .B(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n67), .CI(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n19), .CO(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n18), .S(fu_LIFTING_N654) );
  ADDFX1 fu_LIFTING_mult_96_DP_OP_281_6650_6_U24 ( .A(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n76), .B(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n77), .CI(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n24), .CO(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n23), .S(fu_LIFTING_N649) );
  ADDFX1 fu_LIFTING_mult_96_DP_OP_281_6650_6_U25 ( .A(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n78), .B(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n79), .CI(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n25), .CO(
        fu_LIFTING_mult_96_DP_OP_281_6650_6_n24), .S(fu_LIFTING_N648) );
  EDFFX2 fu_LIFTING_reg_x1_reg_1_ ( .D(n2110), .E(fu_LIFTING_n85), .CK(clk), 
        .Q(fu_LIFTING_reg_x1_1_) );
  EDFFX2 fu_LIFTING_reg_x1_reg_4_ ( .D(n1825), .E(fu_LIFTING_n85), .CK(clk), 
        .Q(fu_LIFTING_reg_x1_4_) );
  EDFFX2 fu_LIFTING_reg_x2_reg_3_ ( .D(rf_RF_t1data_wire[3]), .E(
        fu_LIFTING_n244), .CK(clk), .Q(fu_LIFTING_reg_x2_3_) );
  EDFFX2 fu_LIFTING_reg_x2_reg_4_ ( .D(n1825), .E(fu_LIFTING_n244), .CK(clk), 
        .Q(fu_LIFTING_reg_x2_4_) );
  EDFFX2 fu_LIFTING_reg_x1_reg_0_ ( .D(n2111), .E(fu_LIFTING_n85), .CK(clk), 
        .Q(fu_LIFTING_reg_x1_0_) );
  EDFFX2 fu_LIFTING_reg_x1_reg_2_ ( .D(n1810), .E(fu_LIFTING_n85), .CK(clk), 
        .Q(fu_LIFTING_reg_x1_2_) );
  EDFFX2 fu_LIFTING_reg_x1_reg_3_ ( .D(rf_RF_t1data_wire[3]), .E(
        fu_LIFTING_n85), .CK(clk), .Q(fu_LIFTING_reg_x1_3_) );
  EDFFX2 fu_LIFTING_reg_x1_reg_5_ ( .D(rf_RF_t1data_wire[5]), .E(
        fu_LIFTING_n85), .CK(clk), .Q(fu_LIFTING_reg_x1_5_) );
  EDFFX2 fu_LIFTING_reg_x1_reg_6_ ( .D(n1818), .E(fu_LIFTING_n85), .CK(clk), 
        .Q(fu_LIFTING_reg_x1_6_) );
  EDFFX2 fu_LIFTING_reg_x1_reg_7_ ( .D(n1814), .E(fu_LIFTING_n85), .CK(clk), 
        .Q(fu_LIFTING_reg_x1_7_) );
  EDFFX2 fu_LIFTING_reg_x1_reg_8_ ( .D(rf_RF_t1data_wire[8]), .E(
        fu_LIFTING_n85), .CK(clk), .Q(fu_LIFTING_reg_x1_8_) );
  EDFFX2 fu_LIFTING_reg_x2_reg_1_ ( .D(n2110), .E(fu_LIFTING_n244), .CK(clk), 
        .Q(fu_LIFTING_reg_x2_1_) );
  EDFFX2 fu_LIFTING_reg_x2_reg_2_ ( .D(n1810), .E(fu_LIFTING_n244), .CK(clk), 
        .Q(fu_LIFTING_reg_x2_2_) );
  EDFFX2 fu_LIFTING_reg_x2_reg_5_ ( .D(rf_RF_t1data_wire[5]), .E(
        fu_LIFTING_n244), .CK(clk), .Q(fu_LIFTING_reg_x2_5_) );
  EDFFX2 fu_LIFTING_reg_x2_reg_6_ ( .D(n1818), .E(fu_LIFTING_n244), .CK(clk), 
        .Q(fu_LIFTING_reg_x2_6_) );
  EDFFX2 fu_LIFTING_reg_x2_reg_7_ ( .D(n1814), .E(fu_LIFTING_n244), .CK(clk), 
        .Q(fu_LIFTING_reg_x2_7_) );
  EDFFX2 fu_LIFTING_reg_x2_reg_0_ ( .D(n2111), .E(fu_LIFTING_n244), .CK(clk), 
        .Q(fu_LIFTING_reg_x2_0_) );
  EDFFX2 fu_LIFTING_reg_x1_reg_9_ ( .D(n1812), .E(fu_LIFTING_n85), .CK(clk), 
        .Q(fu_LIFTING_reg_x1_9_) );
  EDFFX2 fu_LIFTING_reg_x1_reg_10_ ( .D(n1816), .E(fu_LIFTING_n85), .CK(clk), 
        .Q(fu_LIFTING_reg_x1_10_) );
  EDFFX2 fu_LIFTING_reg_x1_reg_11_ ( .D(rf_RF_t1data_wire[11]), .E(
        fu_LIFTING_n85), .CK(clk), .Q(fu_LIFTING_reg_x1_11_) );
  EDFFX2 fu_LIFTING_reg_x1_reg_12_ ( .D(n1820), .E(fu_LIFTING_n85), .CK(clk), 
        .Q(fu_LIFTING_reg_x1_12_) );
  EDFFX2 fu_LIFTING_reg_x1_reg_13_ ( .D(n1823), .E(fu_LIFTING_n85), .CK(clk), 
        .Q(fu_LIFTING_reg_x1_13_) );
  EDFFX2 fu_LIFTING_reg_x1_reg_14_ ( .D(rf_RF_t1data_wire[14]), .E(
        fu_LIFTING_n85), .CK(clk), .Q(fu_LIFTING_reg_x1_14_) );
  EDFFX2 fu_LIFTING_reg_x2_reg_8_ ( .D(rf_RF_t1data_wire[8]), .E(
        fu_LIFTING_n244), .CK(clk), .Q(fu_LIFTING_reg_x2_8_) );
  EDFFX2 fu_LIFTING_reg_x2_reg_9_ ( .D(n1812), .E(fu_LIFTING_n244), .CK(clk), 
        .Q(fu_LIFTING_reg_x2_9_) );
  EDFFX2 fu_LIFTING_reg_x2_reg_10_ ( .D(n1816), .E(fu_LIFTING_n244), .CK(clk), 
        .Q(fu_LIFTING_reg_x2_10_) );
  EDFFX2 fu_LIFTING_reg_x2_reg_11_ ( .D(rf_RF_t1data_wire[11]), .E(
        fu_LIFTING_n244), .CK(clk), .Q(fu_LIFTING_reg_x2_11_) );
  EDFFX2 fu_LIFTING_reg_x2_reg_12_ ( .D(n1820), .E(fu_LIFTING_n244), .CK(clk), 
        .Q(fu_LIFTING_reg_x2_12_) );
  EDFFX2 fu_LIFTING_reg_x2_reg_13_ ( .D(n1823), .E(fu_LIFTING_n245), .CK(clk), 
        .Q(fu_LIFTING_reg_x2_13_) );
  EDFFX2 fu_LIFTING_reg_x1_reg_15_ ( .D(rf_RF_t1data_wire[15]), .E(
        fu_LIFTING_n85), .CK(clk), .Q(fu_LIFTING_reg_x1_15_) );
  EDFFX2 fu_LIFTING_reg_x1_reg_16_ ( .D(rf_RF_t1data_wire[16]), .E(
        fu_LIFTING_n85), .CK(clk), .Q(fu_LIFTING_reg_x1_16_) );
  EDFFX2 fu_LIFTING_reg_x1_reg_17_ ( .D(rf_RF_t1data_wire[17]), .E(
        fu_LIFTING_n85), .CK(clk), .Q(fu_LIFTING_reg_x1_17_) );
  EDFFX2 fu_LIFTING_reg_x1_reg_18_ ( .D(rf_RF_t1data_wire[18]), .E(
        fu_LIFTING_n85), .CK(clk), .Q(fu_LIFTING_reg_x1_18_) );
  EDFFX2 fu_LIFTING_reg_x1_reg_19_ ( .D(rf_RF_t1data_wire[19]), .E(
        fu_LIFTING_n85), .CK(clk), .Q(fu_LIFTING_reg_x1_19_) );
  EDFFX2 fu_LIFTING_reg_x1_reg_20_ ( .D(rf_RF_t1data_wire[20]), .E(
        fu_LIFTING_n85), .CK(clk), .Q(fu_LIFTING_reg_x1_20_) );
  EDFFX2 fu_LIFTING_reg_x2_reg_14_ ( .D(rf_RF_t1data_wire[14]), .E(
        fu_LIFTING_n245), .CK(clk), .Q(fu_LIFTING_reg_x2_14_) );
  EDFFX2 fu_LIFTING_reg_x2_reg_15_ ( .D(rf_RF_t1data_wire[15]), .E(
        fu_LIFTING_n245), .CK(clk), .Q(fu_LIFTING_reg_x2_15_) );
  EDFFX2 fu_LIFTING_reg_x2_reg_16_ ( .D(rf_RF_t1data_wire[16]), .E(
        fu_LIFTING_n245), .CK(clk), .Q(fu_LIFTING_reg_x2_16_) );
  EDFFX2 fu_LIFTING_reg_x2_reg_17_ ( .D(rf_RF_t1data_wire[17]), .E(
        fu_LIFTING_n245), .CK(clk), .Q(fu_LIFTING_reg_x2_17_) );
  EDFFX2 fu_LIFTING_reg_x2_reg_18_ ( .D(rf_RF_t1data_wire[18]), .E(
        fu_LIFTING_n245), .CK(clk), .Q(fu_LIFTING_reg_x2_18_) );
  EDFFX2 fu_LIFTING_reg_x2_reg_19_ ( .D(rf_RF_t1data_wire[19]), .E(
        fu_LIFTING_n245), .CK(clk), .Q(fu_LIFTING_reg_x2_19_) );
  EDFFX2 fu_LIFTING_reg_x2_reg_20_ ( .D(rf_RF_t1data_wire[20]), .E(
        fu_LIFTING_n245), .CK(clk), .Q(fu_LIFTING_reg_x2_20_) );
  EDFFX2 fu_LIFTING_reg_x2_reg_21_ ( .D(rf_RF_t1data_wire[21]), .E(
        fu_LIFTING_n245), .CK(clk), .Q(fu_LIFTING_reg_x2_21_) );
  EDFFX2 fu_LIFTING_reg_x1_reg_21_ ( .D(rf_RF_t1data_wire[21]), .E(
        fu_LIFTING_n85), .CK(clk), .Q(fu_LIFTING_reg_x1_21_) );
  EDFFX2 fu_LIFTING_reg_x1_reg_22_ ( .D(rf_RF_t1data_wire[22]), .E(
        fu_LIFTING_n85), .CK(clk), .Q(fu_LIFTING_reg_x1_22_) );
  EDFFX2 fu_LIFTING_reg_x1_reg_23_ ( .D(rf_RF_t1data_wire[23]), .E(
        fu_LIFTING_n85), .CK(clk), .Q(fu_LIFTING_reg_x1_23_) );
  EDFFX2 fu_LIFTING_reg_x1_reg_24_ ( .D(rf_RF_t1data_wire[24]), .E(
        fu_LIFTING_n85), .CK(clk), .Q(fu_LIFTING_reg_x1_24_) );
  EDFFX2 fu_LIFTING_reg_x1_reg_25_ ( .D(rf_RF_t1data_wire[25]), .E(
        fu_LIFTING_n85), .CK(clk), .Q(fu_LIFTING_reg_x1_25_) );
  EDFFX2 fu_LIFTING_reg_x1_reg_26_ ( .D(rf_RF_t1data_wire[26]), .E(
        fu_LIFTING_N961), .CK(clk), .Q(fu_LIFTING_reg_x1_26_) );
  EDFFX2 fu_LIFTING_reg_x1_reg_27_ ( .D(rf_RF_t1data_wire[27]), .E(
        fu_LIFTING_N961), .CK(clk), .Q(fu_LIFTING_reg_x1_27_) );
  EDFFX2 fu_LIFTING_reg_x2_reg_22_ ( .D(rf_RF_t1data_wire[22]), .E(
        fu_LIFTING_n245), .CK(clk), .Q(fu_LIFTING_reg_x2_22_) );
  EDFFX2 fu_LIFTING_reg_x2_reg_23_ ( .D(rf_RF_t1data_wire[23]), .E(
        fu_LIFTING_n245), .CK(clk), .Q(fu_LIFTING_reg_x2_23_) );
  EDFFX2 fu_LIFTING_reg_x2_reg_24_ ( .D(rf_RF_t1data_wire[24]), .E(
        fu_LIFTING_n245), .CK(clk), .Q(fu_LIFTING_reg_x2_24_) );
  EDFFX2 fu_LIFTING_reg_x2_reg_25_ ( .D(rf_RF_t1data_wire[25]), .E(
        fu_LIFTING_n245), .CK(clk), .Q(fu_LIFTING_reg_x2_25_) );
  EDFFX2 fu_LIFTING_reg_x2_reg_26_ ( .D(rf_RF_t1data_wire[26]), .E(
        fu_LIFTING_n244), .CK(clk), .Q(fu_LIFTING_reg_x2_26_) );
  EDFFX2 fu_LIFTING_reg_x2_reg_27_ ( .D(rf_RF_t1data_wire[27]), .E(
        fu_LIFTING_n245), .CK(clk), .Q(fu_LIFTING_reg_x2_27_) );
  EDFFX2 fu_LIFTING_reg_x1_reg_28_ ( .D(rf_RF_t1data_wire[28]), .E(
        fu_LIFTING_n85), .CK(clk), .Q(fu_LIFTING_reg_x1_28_) );
  EDFFX2 fu_LIFTING_reg_x1_reg_29_ ( .D(n1861), .E(fu_LIFTING_n85), .CK(clk), 
        .Q(fu_LIFTING_reg_x1_29_) );
  EDFFX2 fu_LIFTING_reg_x1_reg_30_ ( .D(n1862), .E(fu_LIFTING_n85), .CK(clk), 
        .Q(fu_LIFTING_reg_x1_30_) );
  EDFFX2 fu_LIFTING_reg_x2_reg_28_ ( .D(rf_RF_t1data_wire[28]), .E(
        fu_LIFTING_n244), .CK(clk), .Q(fu_LIFTING_reg_x2_28_) );
  EDFFX2 fu_LIFTING_reg_x2_reg_29_ ( .D(n1861), .E(fu_LIFTING_n245), .CK(clk), 
        .Q(fu_LIFTING_reg_x2_29_) );
  EDFFX2 fu_LIFTING_reg_x2_reg_30_ ( .D(n1862), .E(fu_LIFTING_n244), .CK(clk), 
        .Q(fu_LIFTING_reg_x2_30_) );
  EDFFX2 fu_LIFTING_reg_x2_reg_31_ ( .D(n1860), .E(fu_LIFTING_n245), .CK(clk), 
        .Q(fu_LIFTING_reg_x2_31_) );
  EDFFX2 fu_LIFTING_reg_out_tmp_reg_0_ ( .D(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_0_), .E(fu_LIFTING_n84), .CK(clk), .Q(fu_LIFTING_reg_out_tmp_0_) );
  EDFFX2 fu_LIFTING_reg_out_tmp_reg_1_ ( .D(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_1_), .E(fu_LIFTING_n84), .CK(clk), .Q(fu_LIFTING_reg_out_tmp_1_) );
  EDFFX2 fu_LIFTING_reg_out_tmp_reg_2_ ( .D(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_2_), .E(fu_LIFTING_n84), .CK(clk), .Q(fu_LIFTING_reg_out_tmp_2_) );
  EDFFX2 fu_LIFTING_reg_out_tmp_reg_3_ ( .D(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_3_), .E(fu_LIFTING_n84), .CK(clk), .Q(fu_LIFTING_reg_out_tmp_3_) );
  EDFFX2 fu_LIFTING_reg_out_tmp_reg_4_ ( .D(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_4_), .E(fu_LIFTING_n84), .CK(clk), .Q(fu_LIFTING_reg_out_tmp_4_) );
  EDFFX2 fu_LIFTING_reg_out_tmp_reg_5_ ( .D(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_5_), .E(fu_LIFTING_n84), .CK(clk), .Q(fu_LIFTING_reg_out_tmp_5_) );
  EDFFX2 fu_LIFTING_reg_out_tmp_reg_6_ ( .D(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_6_), .E(fu_LIFTING_n84), .CK(clk), .Q(fu_LIFTING_reg_out_tmp_6_) );
  EDFFX2 fu_LIFTING_reg_out_tmp_reg_7_ ( .D(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_7_), .E(fu_LIFTING_n84), .CK(clk), .Q(fu_LIFTING_reg_out_tmp_7_) );
  EDFFX2 fu_LIFTING_reg_out_tmp_reg_8_ ( .D(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_8_), .E(fu_LIFTING_n84), .CK(clk), .Q(fu_LIFTING_reg_out_tmp_8_) );
  EDFFX2 fu_LIFTING_reg_out_tmp_reg_9_ ( .D(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_9_), .E(fu_LIFTING_n84), .CK(clk), .Q(fu_LIFTING_reg_out_tmp_9_) );
  EDFFX2 fu_LIFTING_reg_out_tmp_reg_10_ ( .D(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_10_), .E(fu_LIFTING_n84), .CK(
        clk), .Q(fu_LIFTING_reg_out_tmp_10_) );
  EDFFX2 fu_LIFTING_reg_out_tmp_reg_11_ ( .D(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_11_), .E(fu_LIFTING_n84), .CK(
        clk), .Q(fu_LIFTING_reg_out_tmp_11_) );
  EDFFX2 fu_LIFTING_reg_out_tmp_reg_12_ ( .D(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_12_), .E(fu_LIFTING_n84), .CK(
        clk), .Q(fu_LIFTING_reg_out_tmp_12_) );
  EDFFX2 fu_LIFTING_reg_out_tmp_reg_13_ ( .D(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_13_), .E(fu_LIFTING_n84), .CK(
        clk), .Q(fu_LIFTING_reg_out_tmp_13_) );
  EDFFX2 fu_LIFTING_reg_out_tmp_reg_14_ ( .D(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_14_), .E(fu_LIFTING_n84), .CK(
        clk), .Q(fu_LIFTING_reg_out_tmp_14_) );
  EDFFX2 fu_LIFTING_reg_out_tmp_reg_15_ ( .D(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_15_), .E(fu_LIFTING_n84), .CK(
        clk), .Q(fu_LIFTING_reg_out_tmp_15_) );
  EDFFX2 fu_LIFTING_reg_out_tmp_reg_16_ ( .D(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_16_), .E(fu_LIFTING_n84), .CK(
        clk), .Q(fu_LIFTING_reg_out_tmp_16_) );
  EDFFX2 fu_LIFTING_reg_out_tmp_reg_17_ ( .D(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_17_), .E(fu_LIFTING_n84), .CK(
        clk), .Q(fu_LIFTING_reg_out_tmp_17_) );
  EDFFX2 fu_LIFTING_reg_out_tmp_reg_18_ ( .D(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_18_), .E(fu_LIFTING_n84), .CK(
        clk), .Q(fu_LIFTING_reg_out_tmp_18_) );
  EDFFX2 fu_LIFTING_reg_out_tmp_reg_19_ ( .D(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_19_), .E(fu_LIFTING_n84), .CK(
        clk), .Q(fu_LIFTING_reg_out_tmp_19_) );
  EDFFX2 fu_LIFTING_reg_out_tmp_reg_20_ ( .D(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_20_), .E(fu_LIFTING_n84), .CK(
        clk), .Q(fu_LIFTING_reg_out_tmp_20_) );
  EDFFX2 fu_LIFTING_reg_out_tmp_reg_21_ ( .D(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_21_), .E(fu_LIFTING_n84), .CK(
        clk), .Q(fu_LIFTING_reg_out_tmp_21_) );
  EDFFX2 fu_LIFTING_reg_out_tmp_reg_22_ ( .D(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_22_), .E(fu_LIFTING_n84), .CK(
        clk), .Q(fu_LIFTING_reg_out_tmp_22_) );
  EDFFX2 fu_LIFTING_reg_out_tmp_reg_23_ ( .D(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_23_), .E(fu_LIFTING_n84), .CK(
        clk), .Q(fu_LIFTING_reg_out_tmp_23_) );
  EDFFX2 fu_LIFTING_reg_out_tmp_reg_24_ ( .D(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_24_), .E(fu_LIFTING_n84), .CK(
        clk), .Q(fu_LIFTING_reg_out_tmp_24_) );
  EDFFX2 fu_LIFTING_reg_out_tmp_reg_25_ ( .D(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_25_), .E(fu_LIFTING_n84), .CK(
        clk), .Q(fu_LIFTING_reg_out_tmp_25_) );
  EDFFX2 fu_LIFTING_reg_out_tmp_reg_26_ ( .D(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_26_), .E(fu_LIFTING_n84), .CK(
        clk), .Q(fu_LIFTING_reg_out_tmp_26_) );
  EDFFX2 fu_LIFTING_reg_out_tmp_reg_27_ ( .D(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_27_), .E(fu_LIFTING_n84), .CK(
        clk), .Q(fu_LIFTING_reg_out_tmp_27_) );
  EDFFX2 fu_LIFTING_reg_out_tmp_reg_28_ ( .D(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_28_), .E(fu_LIFTING_n84), .CK(
        clk), .Q(fu_LIFTING_reg_out_tmp_28_) );
  EDFFX2 fu_LIFTING_reg_out_tmp_reg_29_ ( .D(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_29_), .E(fu_LIFTING_n84), .CK(
        clk), .Q(fu_LIFTING_reg_out_tmp_29_) );
  EDFFX2 fu_LIFTING_reg_out_tmp_reg_30_ ( .D(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_30_), .E(fu_LIFTING_N993), .CK(
        clk), .Q(fu_LIFTING_reg_out_tmp_30_) );
  EDFFX2 fu_LIFTING_reg_x1_reg_31_ ( .D(n1860), .E(fu_LIFTING_n85), .CK(clk), 
        .Q(fu_LIFTING_reg_x1_31_) );
  EDFFX2 fu_LIFTING_reg_out_tmp_reg_31_ ( .D(
        fu_LIFTING_sub_98_DP_OP_282_1544_7_O1_31_), .E(fu_LIFTING_N993), .CK(
        clk), .Q(fu_LIFTING_reg_out_tmp_31_) );
endmodule

